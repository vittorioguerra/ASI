VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

VIA via1_2_1120_340_1_3_300_300
  VIARULE Via1Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal1 via1 metal2 ;
  CUTSPACING 0.08 0.08 ;
  ENCLOSURE 0.035 0.05 0.035 0.035 ;
  ROWCOL 1 3 ;
END via1_2_1120_340_1_3_300_300

VIA via2_3_1120_340_1_3_320_320
  VIARULE Via2Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal2 via2 metal3 ;
  CUTSPACING 0.09 0.09 ;
  ENCLOSURE 0.035 0.035 0.035 0.035 ;
  ROWCOL 1 3 ;
END via2_3_1120_340_1_3_320_320

VIA via3_4_1120_340_1_3_320_320
  VIARULE Via3Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal3 via3 metal4 ;
  CUTSPACING 0.09 0.09 ;
  ENCLOSURE 0.035 0.035 0.035 0.035 ;
  ROWCOL 1 3 ;
END via3_4_1120_340_1_3_320_320

VIA via4_5_1120_340_1_2_600_600
  VIARULE Via4Array-0 ;
  CUTSIZE 0.14 0.14 ;
  LAYERS metal4 via4 metal5 ;
  CUTSPACING 0.16 0.16 ;
  ENCLOSURE 0 0 0 0 ;
  ROWCOL 1 2 ;
END via4_5_1120_340_1_2_600_600

VIA via5_6_1120_340_1_2_600_600
  VIARULE Via5Array-0 ;
  CUTSIZE 0.14 0.14 ;
  LAYERS metal5 via5 metal6 ;
  CUTSPACING 0.16 0.16 ;
  ENCLOSURE 0 0 0.06 0 ;
  ROWCOL 1 2 ;
END via5_6_1120_340_1_2_600_600

MACRO enfasi
  FOREIGN enfasi 0 0 ;
  CLASS BLOCK ;
  SIZE 85 BY 85 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  84.93 31.955 85 32.025 ;
    END
  END clk
  PIN q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 23.835 0.07 23.905 ;
    END
  END q[0]
  PIN q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  60.48 84.93 60.55 85 ;
    END
  END q[10]
  PIN q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  84.93 8.715 85 8.785 ;
    END
  END q[11]
  PIN q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  84.93 78.435 85 78.505 ;
    END
  END q[1]
  PIN q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  13.36 84.93 13.43 85 ;
    END
  END q[2]
  PIN q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 35.595 0.07 35.665 ;
    END
  END q[3]
  PIN q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  76.44 84.93 76.51 85 ;
    END
  END q[4]
  PIN q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 82.075 0.07 82.145 ;
    END
  END q[5]
  PIN q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  47.94 0 48.01 0.07 ;
    END
  END q[6]
  PIN q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 12.355 0.07 12.425 ;
    END
  END q[7]
  PIN q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  79.48 0 79.55 0.07 ;
    END
  END q[8]
  PIN q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  0.82 0 0.89 0.07 ;
    END
  END q[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  16.4 0 16.47 0.07 ;
    END
  END rst
  PIN z[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  28.94 84.93 29.01 85 ;
    END
  END z[0]
  PIN z[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  84.93 20.475 85 20.545 ;
    END
  END z[10]
  PIN z[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  31.98 0 32.05 0.07 ;
    END
  END z[1]
  PIN z[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  84.93 55.195 85 55.265 ;
    END
  END z[2]
  PIN z[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  84.93 66.675 85 66.745 ;
    END
  END z[3]
  PIN z[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 58.835 0.07 58.905 ;
    END
  END z[4]
  PIN z[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  44.9 84.93 44.97 85 ;
    END
  END z[5]
  PIN z[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  63.52 0 63.59 0.07 ;
    END
  END z[6]
  PIN z[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 47.075 0.07 47.145 ;
    END
  END z[7]
  PIN z[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 70.315 0.07 70.385 ;
    END
  END z[8]
  PIN z[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  84.93 43.435 85 43.505 ;
    END
  END z[9]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal6 ;
        RECT  75.29 0 75.85 85 ;
        RECT  65.29 0 65.85 85 ;
        RECT  55.29 0 55.85 85 ;
        RECT  45.29 0 45.85 85 ;
        RECT  35.29 0 35.85 85 ;
        RECT  25.29 0 25.85 85 ;
        RECT  15.29 0 15.85 85 ;
        RECT  5.29 0 5.85 85 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal6 ;
        RECT  80.29 0 80.85 85 ;
        RECT  70.29 0 70.85 85 ;
        RECT  60.29 0 60.85 85 ;
        RECT  50.29 0 50.85 85 ;
        RECT  40.29 0 40.85 85 ;
        RECT  30.29 0 30.85 85 ;
        RECT  20.29 0 20.85 85 ;
        RECT  10.29 0 10.85 85 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
     RECT  0.44 27.195 0.57 27.265 ;
     RECT  0.57 1.315 4.05 84.085 ;
     RECT  4.05 1.015 4.235 84.085 ;
     RECT  4.235 1.155 6.71 84.085 ;
     RECT  6.71 1.155 8.23 84.245 ;
     RECT  8.23 0.035 13.43 84.385 ;
     RECT  13.43 0.035 21.98 84.245 ;
     RECT  21.98 0.035 32.93 84.085 ;
     RECT  32.93 0.035 39.39 84.245 ;
     RECT  39.39 0.035 40.91 84.525 ;
     RECT  40.91 0.035 48.01 84.665 ;
     RECT  48.01 1.015 48.32 84.665 ;
     RECT  48.32 1.015 61.05 84.805 ;
     RECT  61.05 1.015 64.73 84.945 ;
     RECT  64.73 1.015 64.92 84.665 ;
     RECT  64.92 1.155 69.22 84.665 ;
     RECT  69.22 1.155 77.27 84.805 ;
     RECT  77.27 1.315 77.65 84.805 ;
     RECT  77.65 1.315 84.36 84.085 ;
    LAYER metal2 ;
     RECT  63.71 0 63.97 0.035 ;
     RECT  0.82 0.035 0.89 1.015 ;
     RECT  8.23 0.035 8.3 1.015 ;
     RECT  16.4 0.035 16.47 1.015 ;
     RECT  31.98 0.035 32.05 1.015 ;
     RECT  47.94 0.035 48.01 1.015 ;
     RECT  63.52 0.035 63.97 1.015 ;
     RECT  79.48 0.035 79.55 1.155 ;
     RECT  0.82 1.015 4.12 1.33 ;
     RECT  8.23 1.015 19.89 1.33 ;
     RECT  24.57 1.015 24.64 1.33 ;
     RECT  28.56 1.015 32.05 1.33 ;
     RECT  42.05 1.015 42.5 1.33 ;
     RECT  47.94 1.015 52 1.33 ;
     RECT  57.82 1.015 58.27 1.33 ;
     RECT  63.52 1.015 64.92 1.33 ;
     RECT  77.2 1.155 79.55 1.33 ;
     RECT  0.82 1.33 19.89 1.715 ;
     RECT  24.57 1.33 35.8 1.715 ;
     RECT  42.05 1.33 58.27 1.715 ;
     RECT  63.52 1.33 65.8 1.715 ;
     RECT  0.82 1.715 20.65 1.855 ;
     RECT  24.57 1.715 65.8 1.855 ;
     RECT  75.34 1.33 79.55 1.995 ;
     RECT  0.82 1.855 65.8 2.555 ;
     RECT  0.82 2.555 67.77 2.73 ;
     RECT  0.82 2.73 70.8 3.115 ;
     RECT  75.34 1.995 81.83 3.115 ;
     RECT  0.82 3.115 81.83 3.535 ;
     RECT  0.82 3.535 82.78 3.955 ;
     RECT  0.82 3.955 83.54 4.585 ;
     RECT  1.39 4.585 83.54 4.795 ;
     RECT  1.39 4.795 84.11 12.355 ;
     RECT  1.01 12.355 84.11 18.865 ;
     RECT  1.01 18.865 83.35 23.835 ;
     RECT  0.82 23.835 83.35 24.815 ;
     RECT  0.82 24.815 84.11 24.885 ;
     RECT  0.82 24.885 83.92 27.195 ;
     RECT  0.44 27.195 83.92 30.415 ;
     RECT  0.44 30.415 84.11 31.815 ;
     RECT  0.44 31.815 84.49 51.135 ;
     RECT  0.44 51.135 84.68 76.125 ;
     RECT  0.63 76.125 84.68 76.685 ;
     RECT  0.63 76.685 84.11 80.045 ;
     RECT  0.63 80.045 83.73 80.465 ;
     RECT  1.01 80.465 82.78 81.025 ;
     RECT  1.01 81.025 1.08 82.145 ;
     RECT  5.34 81.025 82.78 82.67 ;
     RECT  28.94 82.67 82.78 82.845 ;
     RECT  38.63 82.845 82.78 82.985 ;
     RECT  38.63 82.985 82.02 83.265 ;
     RECT  38.82 83.265 80.8 83.405 ;
     RECT  6.71 82.67 21.98 84.07 ;
     RECT  28.94 82.845 33 84.07 ;
     RECT  39.01 83.405 80.8 84.07 ;
     RECT  6.71 84.07 17.04 84.245 ;
     RECT  21.91 84.07 21.98 84.245 ;
     RECT  32.93 84.07 33 84.245 ;
     RECT  39.01 84.07 77.65 84.245 ;
     RECT  8.23 84.245 8.3 84.385 ;
     RECT  69.22 84.245 77.65 84.385 ;
     RECT  39.39 84.245 40.98 84.525 ;
     RECT  52.88 84.245 64.73 84.525 ;
     RECT  40.91 84.525 40.98 84.665 ;
     RECT  56.49 84.525 64.73 84.665 ;
     RECT  73.78 84.385 77.65 84.665 ;
     RECT  44.9 84.245 48.39 84.805 ;
     RECT  58.39 84.665 64.73 84.805 ;
     RECT  69.22 84.385 69.29 84.805 ;
     RECT  76.44 84.665 77.65 84.805 ;
     RECT  59.15 84.805 64.73 84.945 ;
     RECT  13.36 84.245 13.43 84.965 ;
     RECT  28.94 84.07 29.01 84.965 ;
     RECT  44.9 84.805 44.97 84.965 ;
     RECT  60.48 84.945 60.55 84.965 ;
     RECT  76.44 84.805 76.51 84.965 ;
    LAYER metal3 ;
     RECT  0 58.975 0.035 59.185 ;
     RECT  0.035 82.075 0.63 82.145 ;
     RECT  0.035 35.595 0.82 35.665 ;
     RECT  0.82 53.235 1.01 53.305 ;
     RECT  0.035 58.835 1.01 59.185 ;
     RECT  0.63 80.395 1.08 82.145 ;
     RECT  1.01 15.715 1.2 15.785 ;
     RECT  1.01 20.615 1.2 20.685 ;
     RECT  0.82 35.595 1.2 36.225 ;
     RECT  0.035 47.075 1.2 47.145 ;
     RECT  0.44 76.055 1.2 76.125 ;
     RECT  0.035 12.355 1.39 12.425 ;
     RECT  1.2 15.715 1.39 16.485 ;
     RECT  1.01 53.235 1.39 55.545 ;
     RECT  1.39 15.715 1.58 17.045 ;
     RECT  1.2 20.195 1.58 20.685 ;
     RECT  0.035 23.835 1.58 23.905 ;
     RECT  1.2 35.595 1.58 38.185 ;
     RECT  1.39 41.195 1.58 41.265 ;
     RECT  1.2 46.655 1.58 47.145 ;
     RECT  1.01 58.555 1.58 59.185 ;
     RECT  0.035 70.315 1.58 70.385 ;
     RECT  1.58 41.195 1.77 47.705 ;
     RECT  1.58 70.315 1.77 72.065 ;
     RECT  1.2 76.055 1.77 76.685 ;
     RECT  1.39 7.595 1.96 12.425 ;
     RECT  1.58 15.715 1.96 24.465 ;
     RECT  1.77 41.195 1.96 47.985 ;
     RECT  1.39 50.855 1.96 55.545 ;
     RECT  1.58 58.555 1.96 61.005 ;
     RECT  1.58 34.195 2.15 38.185 ;
     RECT  1.96 41.195 2.15 55.545 ;
     RECT  1.96 58.555 2.15 62.265 ;
     RECT  1.96 7.595 2.34 24.605 ;
     RECT  2.15 29.995 2.34 38.185 ;
     RECT  2.15 41.195 2.34 62.405 ;
     RECT  2.15 66.675 2.34 66.745 ;
     RECT  1.77 70.315 2.34 76.685 ;
     RECT  1.08 80.395 2.34 80.465 ;
     RECT  2.34 7.595 2.53 38.185 ;
     RECT  2.34 41.195 2.53 80.465 ;
     RECT  2.53 7.595 4.43 80.465 ;
     RECT  4.43 7.595 4.81 81.025 ;
     RECT  4.81 7.315 5.34 81.025 ;
     RECT  5.34 1.33 5.8 82.67 ;
     RECT  5.8 3.255 9.18 81.025 ;
     RECT  9.18 2.555 10.34 81.025 ;
     RECT  10.34 2.555 10.51 84.07 ;
     RECT  10.51 1.995 10.8 84.07 ;
     RECT  10.8 1.995 11.34 36.925 ;
     RECT  10.8 39.795 11.34 81.025 ;
     RECT  11.34 2.275 13.93 36.925 ;
     RECT  11.34 39.795 13.93 49.385 ;
     RECT  11.34 52.955 14.31 81.025 ;
     RECT  14.31 52.675 14.69 81.025 ;
     RECT  14.69 52.395 14.88 81.025 ;
     RECT  13.93 2.275 15.26 49.385 ;
     RECT  14.88 52.395 15.26 82.005 ;
     RECT  15.26 2.275 15.34 82.005 ;
     RECT  15.34 1.33 15.8 82.67 ;
     RECT  15.8 2.555 16.28 81.865 ;
     RECT  16.28 2.555 16.65 35.665 ;
     RECT  16.28 38.535 16.65 81.865 ;
     RECT  16.65 2.555 18.87 35.525 ;
     RECT  16.65 38.675 18.87 81.865 ;
     RECT  18.87 1.995 19.63 35.525 ;
     RECT  18.87 38.675 19.63 82.005 ;
     RECT  19.63 1.855 20.2 35.665 ;
     RECT  19.63 38.535 20.2 82.005 ;
     RECT  20.2 1.855 20.34 82.005 ;
     RECT  20.34 1.855 20.8 84.07 ;
     RECT  20.8 1.855 21.41 82.005 ;
     RECT  21.41 1.855 22.17 70.805 ;
     RECT  22.17 1.855 25.14 69.545 ;
     RECT  21.41 73.815 25.14 82.005 ;
     RECT  25.14 1.855 25.34 82.005 ;
     RECT  25.34 1.33 25.8 82.67 ;
     RECT  25.8 1.715 29.51 80.745 ;
     RECT  29.51 1.715 29.96 82.005 ;
     RECT  29.96 1.855 30.34 82.005 ;
     RECT  30.34 1.855 30.8 84.07 ;
     RECT  30.8 1.855 31.29 82.285 ;
     RECT  31.29 2.275 31.86 82.285 ;
     RECT  31.86 3.675 35.34 82.285 ;
     RECT  35.34 1.33 35.8 82.67 ;
     RECT  35.8 1.715 37.11 82.67 ;
     RECT  37.11 1.715 38.82 83.265 ;
     RECT  38.82 1.715 40.34 83.405 ;
     RECT  40.34 1.715 40.8 84.07 ;
     RECT  40.8 1.715 45.34 83.545 ;
     RECT  45.34 1.33 45.8 83.545 ;
     RECT  45.8 1.855 50.34 83.545 ;
     RECT  50.34 1.855 50.8 84.07 ;
     RECT  50.8 1.855 55.34 83.545 ;
     RECT  55.34 1.33 55.8 83.545 ;
     RECT  55.8 1.855 57.51 83.545 ;
     RECT  57.51 1.995 59.15 83.545 ;
     RECT  59.15 1.995 60.55 84.945 ;
     RECT  60.55 1.995 60.8 84.07 ;
     RECT  60.8 1.995 61.94 83.405 ;
     RECT  61.94 1.855 62.76 83.405 ;
     RECT  62.76 1.715 65.11 83.405 ;
     RECT  65.11 1.715 65.34 83.265 ;
     RECT  65.34 1.33 65.68 83.265 ;
     RECT  65.68 1.33 65.8 82.67 ;
     RECT  65.8 3.535 65.87 82.285 ;
     RECT  65.87 4.515 67.01 82.285 ;
     RECT  67.01 4.935 70.34 82.285 ;
     RECT  70.34 2.73 70.8 84.07 ;
     RECT  70.8 4.795 73.78 83.265 ;
     RECT  73.78 4.515 74.8 83.265 ;
     RECT  74.8 4.515 75.34 82.67 ;
     RECT  75.34 1.33 75.8 82.67 ;
     RECT  75.8 4.515 76.13 82.145 ;
     RECT  76.13 4.515 76.32 82.005 ;
     RECT  76.32 4.515 79.67 70.945 ;
     RECT  76.32 74.795 79.67 82.005 ;
     RECT  79.67 4.515 80.34 82.005 ;
     RECT  80.34 2.73 80.8 84.07 ;
     RECT  80.8 4.795 81.26 28.385 ;
     RECT  80.8 31.815 81.26 83.265 ;
     RECT  81.26 4.935 81.83 8.785 ;
     RECT  81.26 12.215 81.83 28.385 ;
     RECT  81.26 31.815 81.83 79.065 ;
     RECT  81.83 7.315 82.02 8.785 ;
     RECT  81.26 83.195 82.02 83.265 ;
     RECT  82.02 7.595 82.21 8.785 ;
     RECT  81.83 25.795 82.21 28.385 ;
     RECT  81.83 31.815 82.21 51.485 ;
     RECT  82.21 40.775 82.4 51.485 ;
     RECT  81.83 55.055 82.4 78.505 ;
     RECT  81.83 12.215 82.59 21.665 ;
     RECT  82.21 25.935 82.59 28.385 ;
     RECT  82.4 58.555 82.59 72.065 ;
     RECT  82.59 12.215 82.78 20.545 ;
     RECT  82.59 25.935 82.78 27.265 ;
     RECT  82.4 40.915 82.78 51.485 ;
     RECT  82.78 15.155 82.97 20.545 ;
     RECT  82.21 31.815 82.97 37.205 ;
     RECT  82.78 41.055 82.97 51.485 ;
     RECT  82.59 65.275 82.97 72.065 ;
     RECT  82.97 41.055 83.16 43.645 ;
     RECT  82.97 66.115 83.16 72.065 ;
     RECT  82.78 12.215 83.35 12.285 ;
     RECT  82.78 26.495 83.35 26.565 ;
     RECT  82.97 47.775 83.35 51.485 ;
     RECT  82.97 17.115 83.54 20.545 ;
     RECT  83.35 47.775 83.54 51.205 ;
     RECT  82.59 58.555 83.54 62.405 ;
     RECT  82.4 77.455 83.54 78.505 ;
     RECT  82.97 31.815 83.73 33.845 ;
     RECT  83.16 66.115 83.73 66.745 ;
     RECT  83.16 70.735 83.73 72.065 ;
     RECT  83.54 59.815 83.92 62.405 ;
     RECT  83.73 66.255 83.92 66.745 ;
     RECT  83.54 17.115 84.11 17.185 ;
     RECT  82.97 37.135 84.3 37.205 ;
     RECT  83.54 47.775 84.3 47.845 ;
     RECT  83.73 31.815 84.49 32.025 ;
     RECT  82.4 55.055 84.49 55.265 ;
     RECT  83.92 62.335 84.49 62.405 ;
     RECT  83.54 51.135 84.68 51.205 ;
     RECT  83.73 70.735 84.68 70.805 ;
     RECT  82.21 8.715 84.965 8.785 ;
     RECT  83.54 20.475 84.965 20.545 ;
     RECT  84.49 31.955 84.965 32.025 ;
     RECT  83.16 43.435 84.965 43.505 ;
     RECT  84.49 55.195 84.965 55.265 ;
     RECT  83.92 66.675 84.965 66.745 ;
     RECT  83.54 78.435 84.965 78.505 ;
    LAYER metal4 ;
     RECT  5.34 1.33 5.8 2.73 ;
     RECT  15.34 1.33 15.8 2.73 ;
     RECT  25.34 1.33 25.8 2.73 ;
     RECT  35.34 1.33 35.8 2.73 ;
     RECT  45.34 1.33 45.8 2.73 ;
     RECT  55.34 1.33 55.8 2.73 ;
     RECT  65.34 1.33 65.8 2.73 ;
     RECT  75.34 1.33 75.8 2.73 ;
     RECT  5.34 2.73 80.8 11.62 ;
     RECT  3.105 11.62 80.8 15.4 ;
     RECT  4.225 15.4 80.8 17.92 ;
     RECT  5.34 17.92 80.8 23.94 ;
     RECT  3.945 23.94 80.8 33.18 ;
     RECT  4.225 33.18 80.8 36.26 ;
     RECT  4.785 36.26 80.8 37.1 ;
     RECT  4.785 37.1 82.485 42.84 ;
     RECT  4.785 42.84 81.645 43.54 ;
     RECT  4.785 43.54 80.8 45.92 ;
     RECT  4.505 45.92 80.8 47.88 ;
     RECT  2.545 47.88 80.8 53.48 ;
     RECT  2.545 53.48 81.645 56.56 ;
     RECT  2.265 56.56 81.645 57.96 ;
     RECT  2.265 57.96 82.205 61.18 ;
     RECT  4.505 61.18 82.205 61.74 ;
     RECT  4.505 61.74 80.8 65.38 ;
     RECT  5.34 65.38 80.8 82.67 ;
     RECT  10.34 82.67 10.8 84.07 ;
     RECT  20.34 82.67 20.8 84.07 ;
     RECT  30.34 82.67 30.8 84.07 ;
     RECT  40.34 82.67 40.8 84.07 ;
     RECT  50.34 82.67 50.8 84.07 ;
     RECT  60.34 82.67 60.8 84.07 ;
     RECT  70.34 82.67 70.8 84.07 ;
     RECT  80.34 82.67 80.8 84.07 ;
    LAYER metal5 ;
     RECT  5.35 1.33 5.79 82.67 ;
     RECT  5.79 2.73 10.35 82.67 ;
     RECT  10.35 2.73 10.79 84.07 ;
     RECT  10.79 2.73 15.35 82.67 ;
     RECT  15.35 1.33 15.79 82.67 ;
     RECT  15.79 2.73 20.35 82.67 ;
     RECT  20.35 2.73 20.79 84.07 ;
     RECT  20.79 2.73 25.35 82.67 ;
     RECT  25.35 1.33 25.79 82.67 ;
     RECT  25.79 2.73 30.35 82.67 ;
     RECT  30.35 2.73 30.79 84.07 ;
     RECT  30.79 2.73 35.35 82.67 ;
     RECT  35.35 1.33 35.79 82.67 ;
     RECT  35.79 2.73 40.35 82.67 ;
     RECT  40.35 2.73 40.79 84.07 ;
     RECT  40.79 2.73 45.35 82.67 ;
     RECT  45.35 1.33 45.79 82.67 ;
     RECT  45.79 2.73 50.35 82.67 ;
     RECT  50.35 2.73 50.79 84.07 ;
     RECT  50.79 2.73 55.35 82.67 ;
     RECT  55.35 1.33 55.79 82.67 ;
     RECT  55.79 2.73 60.35 82.67 ;
     RECT  60.35 2.73 60.79 84.07 ;
     RECT  60.79 2.73 65.35 82.67 ;
     RECT  65.35 1.33 65.79 82.67 ;
     RECT  65.79 2.73 70.35 82.67 ;
     RECT  70.35 2.73 70.79 84.07 ;
     RECT  70.79 2.73 75.35 82.67 ;
     RECT  75.35 1.33 75.79 82.67 ;
     RECT  75.79 2.73 80.35 82.67 ;
     RECT  80.35 2.73 80.79 84.07 ;
    LAYER metal6 ;
     RECT  5.29 0 80.85 85 ;
  END
END enfasi
END LIBRARY
