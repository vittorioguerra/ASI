VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

VIA via1_2_1120_340_1_3_300_300
  VIARULE Via1Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal1 via1 metal2 ;
  CUTSPACING 0.08 0.08 ;
  ENCLOSURE 0.035 0.05 0.035 0.035 ;
  ROWCOL 1 3 ;
END via1_2_1120_340_1_3_300_300

VIA via2_3_1120_340_1_3_320_320
  VIARULE Via2Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal2 via2 metal3 ;
  CUTSPACING 0.09 0.09 ;
  ENCLOSURE 0.035 0.035 0.035 0.035 ;
  ROWCOL 1 3 ;
END via2_3_1120_340_1_3_320_320

VIA via3_4_1120_340_1_3_320_320
  VIARULE Via3Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal3 via3 metal4 ;
  CUTSPACING 0.09 0.09 ;
  ENCLOSURE 0.035 0.035 0.035 0.035 ;
  ROWCOL 1 3 ;
END via3_4_1120_340_1_3_320_320

VIA via4_5_1120_340_1_2_600_600
  VIARULE Via4Array-0 ;
  CUTSIZE 0.14 0.14 ;
  LAYERS metal4 via4 metal5 ;
  CUTSPACING 0.16 0.16 ;
  ENCLOSURE 0 0 0 0 ;
  ROWCOL 1 2 ;
END via4_5_1120_340_1_2_600_600

VIA via5_6_1120_340_1_2_600_600
  VIARULE Via5Array-0 ;
  CUTSIZE 0.14 0.14 ;
  LAYERS metal5 via5 metal6 ;
  CUTSPACING 0.16 0.16 ;
  ENCLOSURE 0 0 0.06 0 ;
  ROWCOL 1 2 ;
END via5_6_1120_340_1_2_600_600

MACRO iir
  FOREIGN iir 0 0 ;
  CLASS BLOCK ;
  SIZE 75 BY 75 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  59.72 74.93 59.79 75 ;
    END
  END clk
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 21.875 0.07 21.945 ;
    END
  END rst
  PIN x[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  16.4 74.93 16.47 75 ;
    END
  END x[0]
  PIN x[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  74.93 63.595 75 63.665 ;
    END
  END x[10]
  PIN x[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  74.93 42.315 75 42.385 ;
    END
  END x[1]
  PIN x[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  74.93 21.035 75 21.105 ;
    END
  END x[2]
  PIN x[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  74.16 74.93 74.23 75 ;
    END
  END x[3]
  PIN x[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  58.58 0 58.65 0.07 ;
    END
  END x[4]
  PIN x[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 32.515 0.07 32.585 ;
    END
  END x[5]
  PIN x[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 11.235 0.07 11.305 ;
    END
  END x[6]
  PIN x[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  73.02 0 73.09 0.07 ;
    END
  END x[7]
  PIN x[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  0.82 0 0.89 0.07 ;
    END
  END x[8]
  PIN x[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  15.26 0 15.33 0.07 ;
    END
  END x[9]
  PIN z[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  30.84 74.93 30.91 75 ;
    END
  END z[0]
  PIN z[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  74.93 10.395 75 10.465 ;
    END
  END z[10]
  PIN z[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  29.7 0 29.77 0.07 ;
    END
  END z[1]
  PIN z[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  1.96 74.93 2.03 75 ;
    END
  END z[2]
  PIN z[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  74.93 52.955 75 53.025 ;
    END
  END z[3]
  PIN z[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 53.795 0.07 53.865 ;
    END
  END z[4]
  PIN z[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  45.28 74.93 45.35 75 ;
    END
  END z[5]
  PIN z[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  44.14 0 44.21 0.07 ;
    END
  END z[6]
  PIN z[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 43.155 0.07 43.225 ;
    END
  END z[7]
  PIN z[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 64.435 0.07 64.505 ;
    END
  END z[8]
  PIN z[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  74.93 31.675 75 31.745 ;
    END
  END z[9]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal6 ;
        RECT  65.29 74.86 65.85 75 ;
        RECT  65.29 0 65.85 0.14 ;
        RECT  55.29 74.86 55.85 75 ;
        RECT  55.29 0 55.85 0.14 ;
        RECT  45.29 74.86 45.85 75 ;
        RECT  45.29 0 45.85 0.14 ;
        RECT  35.29 74.86 35.85 75 ;
        RECT  35.29 0 35.85 0.14 ;
        RECT  25.29 74.86 25.85 75 ;
        RECT  25.29 0 25.85 0.14 ;
        RECT  15.29 74.86 15.85 75 ;
        RECT  15.29 0 15.85 0.14 ;
        RECT  5.29 74.86 5.85 75 ;
        RECT  5.29 0 5.85 0.14 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal6 ;
        RECT  70.29 74.86 70.85 75 ;
        RECT  70.29 0 70.85 0.14 ;
        RECT  60.29 74.86 60.85 75 ;
        RECT  60.29 0 60.85 0.14 ;
        RECT  50.29 74.86 50.85 75 ;
        RECT  50.29 0 50.85 0.14 ;
        RECT  40.29 74.86 40.85 75 ;
        RECT  40.29 0 40.85 0.14 ;
        RECT  30.29 74.86 30.85 75 ;
        RECT  30.29 0 30.85 0.14 ;
        RECT  20.29 74.86 20.85 75 ;
        RECT  20.29 0 20.85 0.14 ;
        RECT  10.29 74.86 10.85 75 ;
        RECT  10.29 0 10.85 0.14 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
     RECT  0.57 1.315 0.82 74.285 ;
     RECT  0.82 1.155 6.33 74.285 ;
     RECT  6.33 0.735 8.23 74.285 ;
     RECT  8.23 0.735 8.8 74.585 ;
     RECT  8.8 0.735 11.08 74.725 ;
     RECT  11.08 0.595 19.82 74.725 ;
     RECT  19.82 0.595 32.43 74.865 ;
     RECT  32.43 0.735 37.18 74.865 ;
     RECT  37.18 0.735 43.45 74.725 ;
     RECT  43.45 1.155 45.35 74.725 ;
     RECT  45.35 1.155 46.8 74.585 ;
     RECT  46.8 0.735 51.17 74.585 ;
     RECT  51.17 0.595 55.23 74.585 ;
     RECT  55.23 0.595 57.32 74.285 ;
     RECT  57.32 1.015 68.15 74.285 ;
     RECT  68.15 1.315 74.48 74.285 ;
     RECT  74.48 14.595 74.61 14.665 ;
    LAYER metal2 ;
     RECT  72.07 0 72.9 0.035 ;
     RECT  72.07 0.035 73.09 0.245 ;
     RECT  29.7 0.035 29.77 0.595 ;
     RECT  58.58 0.035 58.65 0.595 ;
     RECT  44.14 0.035 44.21 0.735 ;
     RECT  51.17 0.595 51.24 0.735 ;
     RECT  57.25 0.595 58.65 0.735 ;
     RECT  11.08 0.595 11.15 0.875 ;
     RECT  43.38 0.735 46.87 0.875 ;
     RECT  56.11 0.735 58.65 0.875 ;
     RECT  10.89 0.875 11.15 1.015 ;
     RECT  15.26 0.035 15.33 1.015 ;
     RECT  43.38 0.875 47.25 1.015 ;
     RECT  51.17 0.735 51.43 1.015 ;
     RECT  55.92 0.875 58.65 1.015 ;
     RECT  6.33 0.735 6.4 1.155 ;
     RECT  10.89 1.015 15.33 1.155 ;
     RECT  28.94 0.595 32.43 1.155 ;
     RECT  43.38 1.015 51.43 1.155 ;
     RECT  55.92 1.015 61.12 1.155 ;
     RECT  68.08 1.015 68.15 1.155 ;
     RECT  0.82 0.035 0.89 1.225 ;
     RECT  6.33 1.155 19.13 1.33 ;
     RECT  23.62 1.155 34.71 1.33 ;
     RECT  5.34 1.33 19.13 1.715 ;
     RECT  23.62 1.33 35.8 1.715 ;
     RECT  5.34 1.715 38.7 1.995 ;
     RECT  43.38 1.155 68.15 1.995 ;
     RECT  72.07 0.245 72.33 1.995 ;
     RECT  4.24 1.995 72.33 4.095 ;
     RECT  4.24 4.095 72.71 4.795 ;
     RECT  4.24 4.795 73.28 4.865 ;
     RECT  4.24 4.865 73.09 9.135 ;
     RECT  2.34 9.135 73.47 10.395 ;
     RECT  2.15 10.395 74.42 10.675 ;
     RECT  1.96 10.675 74.42 14.595 ;
     RECT  1.58 14.595 74.61 14.805 ;
     RECT  2.34 14.805 74.61 18.795 ;
     RECT  2.15 18.795 74.61 21.105 ;
     RECT  2.15 21.105 74.42 22.855 ;
     RECT  1.96 22.855 74.42 23.485 ;
     RECT  2.15 23.485 74.42 27.055 ;
     RECT  2.15 27.055 74.61 31.675 ;
     RECT  2.15 31.675 74.99 35.315 ;
     RECT  1.96 35.315 74.99 35.595 ;
     RECT  1.77 35.595 74.99 36.715 ;
     RECT  1.58 36.715 74.99 36.855 ;
     RECT  1.2 36.855 74.99 37.275 ;
     RECT  1.01 37.275 74.99 40.845 ;
     RECT  1.77 40.845 74.99 45.115 ;
     RECT  1.58 45.115 74.99 48.335 ;
     RECT  1.58 48.335 74.8 49.595 ;
     RECT  1.39 49.595 74.8 49.665 ;
     RECT  1.58 49.665 74.8 53.865 ;
     RECT  1.58 53.865 74.42 56.245 ;
     RECT  1.58 56.245 72.71 58.135 ;
     RECT  1.01 58.135 72.71 59.045 ;
     RECT  1.39 59.045 72.71 62.335 ;
     RECT  1.39 62.335 73.09 62.825 ;
     RECT  1.58 62.825 73.09 63.665 ;
     RECT  1.96 63.665 73.09 69.265 ;
     RECT  1.96 69.265 65.87 69.545 ;
     RECT  70.34 69.265 73.09 72.87 ;
     RECT  71.5 72.87 73.09 73.395 ;
     RECT  71.5 73.395 74.23 73.465 ;
     RECT  1.96 69.545 65.8 73.745 ;
     RECT  1.96 73.745 48.39 73.885 ;
     RECT  59.72 73.745 65.8 73.885 ;
     RECT  29.7 73.885 48.39 74.025 ;
     RECT  1.96 73.885 25.8 74.27 ;
     RECT  53.07 73.745 55.8 74.27 ;
     RECT  65.34 73.885 65.8 74.27 ;
     RECT  8.23 74.27 23.5 74.445 ;
     RECT  29.7 74.025 47.82 74.445 ;
     RECT  53.07 74.27 55.23 74.445 ;
     RECT  8.23 74.445 10.01 74.585 ;
     RECT  14.31 74.445 23.5 74.585 ;
     RECT  35.02 74.445 45.35 74.585 ;
     RECT  55.16 74.445 55.23 74.585 ;
     RECT  8.8 74.585 8.87 74.725 ;
     RECT  16.4 74.585 23.5 74.725 ;
     RECT  35.02 74.585 40.22 74.725 ;
     RECT  16.4 74.725 19.89 74.865 ;
     RECT  29.7 74.445 30.91 74.865 ;
     RECT  37.11 74.725 37.18 74.865 ;
     RECT  1.96 74.27 2.03 74.965 ;
     RECT  16.4 74.865 16.47 74.965 ;
     RECT  30.84 74.865 30.91 74.965 ;
     RECT  45.28 74.585 45.35 74.965 ;
     RECT  59.72 73.885 59.79 74.965 ;
     RECT  74.16 73.465 74.23 74.965 ;
    LAYER metal3 ;
     RECT  0 21.315 0.035 21.805 ;
     RECT  0 64.155 0.035 64.365 ;
     RECT  0.035 43.155 1.01 43.225 ;
     RECT  1.01 58.135 1.39 58.205 ;
     RECT  0.035 53.795 1.58 53.865 ;
     RECT  1.39 58.135 1.58 59.465 ;
     RECT  1.01 37.975 1.77 43.225 ;
     RECT  0.035 11.235 1.96 11.305 ;
     RECT  0.035 21.315 1.96 21.945 ;
     RECT  0.035 64.155 1.96 64.505 ;
     RECT  1.96 10.395 2.03 11.305 ;
     RECT  1.58 53.795 2.15 54.845 ;
     RECT  1.58 58.135 2.15 59.885 ;
     RECT  1.58 14.595 2.34 14.665 ;
     RECT  0.035 32.515 2.34 32.585 ;
     RECT  1.77 35.595 2.34 43.225 ;
     RECT  2.15 53.795 2.34 59.885 ;
     RECT  1.96 62.755 2.34 64.505 ;
     RECT  2.34 14.455 2.53 14.665 ;
     RECT  2.34 53.795 2.72 64.505 ;
     RECT  2.03 10.395 3.1 10.465 ;
     RECT  2.34 32.375 3.1 32.585 ;
     RECT  2.72 53.795 3.1 65.065 ;
     RECT  3.1 31.535 3.29 32.585 ;
     RECT  2.34 35.595 3.29 46.865 ;
     RECT  3.1 53.795 3.29 65.345 ;
     RECT  3.29 53.795 3.48 66.605 ;
     RECT  3.29 31.535 3.67 46.865 ;
     RECT  3.48 52.115 3.67 66.605 ;
     RECT  3.67 31.535 4.05 66.605 ;
     RECT  2.53 14.175 4.24 14.665 ;
     RECT  1.96 18.795 4.24 21.945 ;
     RECT  4.05 29.155 4.24 66.605 ;
     RECT  4.24 29.155 4.43 69.265 ;
     RECT  3.1 9.135 4.62 10.465 ;
     RECT  4.24 14.175 4.62 21.945 ;
     RECT  4.43 28.735 4.62 69.265 ;
     RECT  4.62 8.715 4.81 10.465 ;
     RECT  4.81 7.595 5 10.465 ;
     RECT  4.62 13.895 5 21.945 ;
     RECT  5 7.595 5.34 24.325 ;
     RECT  4.62 27.195 5.34 69.405 ;
     RECT  5.34 1.33 5.8 74.27 ;
     RECT  5.8 1.995 8.61 73.605 ;
     RECT  8.61 1.995 8.68 73.885 ;
     RECT  8.68 2.73 9.25 73.885 ;
     RECT  9.25 2.73 9.82 73.605 ;
     RECT  9.82 2.73 10.8 72.87 ;
     RECT  10.8 3.395 14.31 70.805 ;
     RECT  14.31 3.395 14.88 71.785 ;
     RECT  14.88 3.395 15.34 73.325 ;
     RECT  15.34 1.33 15.8 74.27 ;
     RECT  15.8 3.115 16.47 73.605 ;
     RECT  16.47 3.115 18.37 73.465 ;
     RECT  18.37 3.115 20.34 73.325 ;
     RECT  20.34 2.73 20.8 73.325 ;
     RECT  20.8 3.115 22.86 73.325 ;
     RECT  22.86 3.115 24.57 73.885 ;
     RECT  24.57 2.135 25.34 73.885 ;
     RECT  25.34 1.33 25.8 74.27 ;
     RECT  25.8 1.855 28.44 73.605 ;
     RECT  28.44 1.855 28.82 73.325 ;
     RECT  28.82 1.855 30.8 72.87 ;
     RECT  30.8 1.855 30.91 72.345 ;
     RECT  30.91 1.855 31.86 71.925 ;
     RECT  31.86 1.995 35.34 71.925 ;
     RECT  35.34 1.33 35.8 74.27 ;
     RECT  35.8 1.995 37.18 72.065 ;
     RECT  37.18 2.135 40.34 72.065 ;
     RECT  40.34 2.135 40.91 72.87 ;
     RECT  40.91 2.135 41.67 73.605 ;
     RECT  41.67 1.995 42.24 73.605 ;
     RECT  42.24 1.995 43.76 73.885 ;
     RECT  43.76 1.855 45.34 73.885 ;
     RECT  45.34 1.33 45.8 74.27 ;
     RECT  45.8 1.995 48.39 74.025 ;
     RECT  48.39 1.995 50.41 73.605 ;
     RECT  50.41 1.855 55.34 73.605 ;
     RECT  55.34 1.33 55.8 74.27 ;
     RECT  55.8 1.995 55.99 73.605 ;
     RECT  55.99 1.995 56.75 73.465 ;
     RECT  56.75 1.995 57.51 72.625 ;
     RECT  57.51 2.975 60.34 72.625 ;
     RECT  60.34 2.73 61.43 72.87 ;
     RECT  61.43 2.73 62.45 73.605 ;
     RECT  62.45 2.73 63.14 46.725 ;
     RECT  63.14 1.715 65.34 46.725 ;
     RECT  62.45 49.595 65.34 73.605 ;
     RECT  65.34 1.33 65.8 74.27 ;
     RECT  65.8 3.395 70.34 69.265 ;
     RECT  70.34 2.73 70.8 72.87 ;
     RECT  70.8 3.395 70.81 12.005 ;
     RECT  70.81 3.395 71.38 11.025 ;
     RECT  70.8 14.875 71.38 63.665 ;
     RECT  71.38 57.715 71.76 58.065 ;
     RECT  71.38 3.395 71.95 10.605 ;
     RECT  71.76 57.995 71.95 58.065 ;
     RECT  71.38 14.875 72.14 54.285 ;
     RECT  71.95 3.395 72.33 6.405 ;
     RECT  71.95 10.395 72.33 10.605 ;
     RECT  72.14 14.875 72.33 34.545 ;
     RECT  72.33 4.655 72.52 6.405 ;
     RECT  72.14 38.535 72.52 44.625 ;
     RECT  70.8 71.995 72.52 72.065 ;
     RECT  72.52 40.075 72.71 44.625 ;
     RECT  72.33 14.875 72.9 21.665 ;
     RECT  72.52 6.335 73.09 6.405 ;
     RECT  72.33 25.935 73.28 34.545 ;
     RECT  72.71 41.195 73.28 44.625 ;
     RECT  72.14 48.475 73.28 54.285 ;
     RECT  73.28 41.195 73.47 43.925 ;
     RECT  72.9 17.535 73.66 21.665 ;
     RECT  73.28 25.935 73.66 28.805 ;
     RECT  73.28 31.675 73.66 34.545 ;
     RECT  73.66 18.655 73.85 21.665 ;
     RECT  73.28 50.855 73.85 54.285 ;
     RECT  73.85 20.195 74.04 21.665 ;
     RECT  73.66 31.675 74.04 33.145 ;
     RECT  73.85 51.415 74.04 53.865 ;
     RECT  74.04 20.195 74.23 21.105 ;
     RECT  73.66 27.055 74.61 27.125 ;
     RECT  73.47 41.195 74.61 42.385 ;
     RECT  74.04 52.955 74.8 53.865 ;
     RECT  72.33 10.395 74.965 10.465 ;
     RECT  74.23 21.035 74.965 21.105 ;
     RECT  74.04 31.675 74.965 31.745 ;
     RECT  74.61 42.315 74.965 42.385 ;
     RECT  74.8 52.955 74.965 53.725 ;
     RECT  71.38 63.595 74.965 63.665 ;
     RECT  74.965 53.095 75 53.725 ;
    LAYER metal4 ;
     RECT  45.34 1.33 45.8 2.24 ;
     RECT  5.34 1.33 5.8 2.73 ;
     RECT  15.34 1.33 15.8 2.73 ;
     RECT  25.34 1.33 25.8 2.73 ;
     RECT  35.34 1.33 35.8 2.73 ;
     RECT  42.025 2.24 45.8 2.73 ;
     RECT  55.34 1.33 55.8 2.73 ;
     RECT  65.34 1.33 65.8 2.73 ;
     RECT  5.34 2.73 70.8 57.68 ;
     RECT  3.665 57.68 70.8 58.94 ;
     RECT  3.385 58.94 70.8 60.9 ;
     RECT  5.34 60.9 70.8 72.87 ;
     RECT  15.34 72.87 16.405 73.64 ;
     RECT  5.34 72.87 5.8 74.27 ;
     RECT  15.34 73.64 15.8 74.27 ;
     RECT  25.34 72.87 25.8 74.27 ;
     RECT  35.34 72.87 35.8 74.27 ;
     RECT  45.34 72.87 45.8 74.27 ;
     RECT  55.34 72.87 55.8 74.27 ;
     RECT  65.34 72.87 65.8 74.27 ;
    LAYER metal5 ;
     RECT  5.35 1.33 5.79 74.27 ;
     RECT  5.79 2.73 15.35 72.87 ;
     RECT  15.35 1.33 15.79 74.27 ;
     RECT  15.79 2.73 25.35 72.87 ;
     RECT  25.35 1.33 25.79 74.27 ;
     RECT  25.79 2.73 35.35 72.87 ;
     RECT  35.35 1.33 35.79 74.27 ;
     RECT  35.79 2.73 45.35 72.87 ;
     RECT  45.35 1.33 45.79 74.27 ;
     RECT  45.79 2.73 55.35 72.87 ;
     RECT  55.35 1.33 55.79 74.27 ;
     RECT  55.79 2.73 65.35 72.87 ;
     RECT  65.35 1.33 65.79 74.27 ;
     RECT  65.79 2.73 70.79 72.87 ;
    LAYER metal6 ;
     RECT  5.29 0 70.85 75 ;
  END
END iir
END LIBRARY
