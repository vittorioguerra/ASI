module iir (clk,
    rst,
    x,
    z);
 input clk;
 input rst;
 input [10:0] x;
 output [10:0] z;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire \coll_reg[0] ;
 wire \coll_reg[10] ;
 wire \coll_reg[1] ;
 wire \coll_reg[2] ;
 wire \coll_reg[3] ;
 wire \coll_reg[4] ;
 wire \coll_reg[5] ;
 wire \coll_reg[6] ;
 wire \coll_reg[7] ;
 wire \coll_reg[8] ;
 wire \coll_reg[9] ;
 wire \in_reg1[0] ;
 wire \in_reg1[10] ;
 wire \in_reg1[1] ;
 wire \in_reg1[2] ;
 wire \in_reg1[3] ;
 wire \in_reg1[4] ;
 wire \in_reg1[5] ;
 wire \in_reg1[6] ;
 wire \in_reg1[7] ;
 wire \in_reg1[8] ;
 wire \in_reg1[9] ;
 wire \section_1.t1[0] ;
 wire \section_1.t1[1] ;
 wire \section_1.t1[2] ;
 wire \section_1.t1[3] ;
 wire \section_1.t1[4] ;
 wire \section_1.xn1[10] ;
 wire \section_1.xn1[5] ;
 wire \section_1.xn1[6] ;
 wire \section_1.xn1[7] ;
 wire \section_1.xn1[8] ;
 wire \section_1.xn1[9] ;
 wire \section_1.xn2[0] ;
 wire \section_1.xn2[10] ;
 wire \section_1.xn2[1] ;
 wire \section_1.xn2[2] ;
 wire \section_1.xn2[3] ;
 wire \section_1.xn2[4] ;
 wire \section_1.xn2[5] ;
 wire \section_1.xn2[6] ;
 wire \section_1.xn2[7] ;
 wire \section_1.xn2[8] ;
 wire \section_1.xn2[9] ;
 wire \section_1.yn2[0] ;
 wire \section_1.yn2[10] ;
 wire \section_1.yn2[1] ;
 wire \section_1.yn2[2] ;
 wire \section_1.yn2[3] ;
 wire \section_1.yn2[4] ;
 wire \section_1.yn2[5] ;
 wire \section_1.yn2[6] ;
 wire \section_1.yn2[7] ;
 wire \section_1.yn2[8] ;
 wire \section_1.yn2[9] ;
 wire \section_2.xn2[0] ;
 wire \section_2.xn2[10] ;
 wire \section_2.xn2[1] ;
 wire \section_2.xn2[2] ;
 wire \section_2.xn2[3] ;
 wire \section_2.xn2[4] ;
 wire \section_2.xn2[5] ;
 wire \section_2.xn2[6] ;
 wire \section_2.xn2[7] ;
 wire \section_2.xn2[8] ;
 wire \section_2.xn2[9] ;
 wire \section_2.yn2[0] ;
 wire \section_2.yn2[10] ;
 wire \section_2.yn2[1] ;
 wire \section_2.yn2[2] ;
 wire \section_2.yn2[3] ;
 wire \section_2.yn2[4] ;
 wire \section_2.yn2[5] ;
 wire \section_2.yn2[6] ;
 wire \section_2.yn2[7] ;
 wire \section_2.yn2[8] ;
 wire \section_2.yn2[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;

 INV_X1 _3015_ (.A(rst),
    .ZN(_1253_));
 XOR2_X1 _3016_ (.A(\section_2.yn2[10] ),
    .B(\section_2.yn2[8] ),
    .Z(_1264_));
 XNOR2_X1 _3017_ (.A(z[1]),
    .B(z[0]),
    .ZN(_1275_));
 INV_X1 _3018_ (.A(net91),
    .ZN(_1286_));
 NOR3_X1 _3019_ (.A1(\coll_reg[2] ),
    .A2(\coll_reg[1] ),
    .A3(\coll_reg[0] ),
    .ZN(_1297_));
 XNOR2_X1 _3020_ (.A(_1286_),
    .B(_1297_),
    .ZN(_1308_));
 XNOR2_X1 _3021_ (.A(\section_1.yn2[2] ),
    .B(_1308_),
    .ZN(_1319_));
 INV_X1 _3022_ (.A(net82),
    .ZN(_1330_));
 NAND2_X1 _3023_ (.A1(\coll_reg[2] ),
    .A2(\coll_reg[1] ),
    .ZN(_1341_));
 XOR2_X1 _3024_ (.A(\coll_reg[2] ),
    .B(\coll_reg[0] ),
    .Z(_1352_));
 OR2_X1 _3025_ (.A1(\coll_reg[1] ),
    .A2(_1352_),
    .ZN(_1363_));
 NAND2_X1 _3026_ (.A1(_1341_),
    .A2(_1363_),
    .ZN(_1374_));
 XOR2_X1 _3027_ (.A(\coll_reg[1] ),
    .B(\coll_reg[0] ),
    .Z(_1385_));
 NAND2_X1 _3028_ (.A1(\section_1.yn2[0] ),
    .A2(_1385_),
    .ZN(_1396_));
 XNOR2_X1 _3029_ (.A(_1330_),
    .B(_1374_),
    .ZN(_1407_));
 OAI22_X1 _3030_ (.A1(_1330_),
    .A2(_1374_),
    .B1(_1396_),
    .B2(_1407_),
    .ZN(_1418_));
 XNOR2_X1 _3031_ (.A(_1319_),
    .B(_1418_),
    .ZN(_1429_));
 INV_X1 _3032_ (.A(\section_2.xn2[3] ),
    .ZN(_1440_));
 XNOR2_X1 _3033_ (.A(_1440_),
    .B(_1429_),
    .ZN(_1451_));
 INV_X1 _3034_ (.A(\section_2.xn2[2] ),
    .ZN(_1462_));
 OAI22_X1 _3035_ (.A1(_0021_),
    .A2(_1429_),
    .B1(_1451_),
    .B2(_1462_),
    .ZN(_1473_));
 INV_X1 _3036_ (.A(\section_2.xn2[4] ),
    .ZN(_1484_));
 NOR2_X1 _3037_ (.A1(_1396_),
    .A2(_1407_),
    .ZN(_1495_));
 NAND2_X1 _3038_ (.A1(_1319_),
    .A2(_1495_),
    .ZN(_1506_));
 NAND4_X1 _3039_ (.A1(\section_1.yn2[1] ),
    .A2(_1341_),
    .A3(_1319_),
    .A4(_1363_),
    .ZN(_1517_));
 INV_X1 _3040_ (.A(net71),
    .ZN(_1528_));
 OR2_X1 _3041_ (.A1(_1528_),
    .A2(_1308_),
    .ZN(_1539_));
 INV_X1 _3042_ (.A(net116),
    .ZN(_1550_));
 NAND2_X1 _3043_ (.A1(\coll_reg[3] ),
    .A2(\coll_reg[2] ),
    .ZN(_1561_));
 NOR2_X1 _3044_ (.A1(_1550_),
    .A2(_1561_),
    .ZN(_1572_));
 NAND2_X1 _3045_ (.A1(\coll_reg[0] ),
    .A2(_1572_),
    .ZN(_1583_));
 XOR2_X1 _3046_ (.A(\coll_reg[4] ),
    .B(\coll_reg[3] ),
    .Z(_1594_));
 XNOR2_X1 _3047_ (.A(\coll_reg[2] ),
    .B(_1594_),
    .ZN(_1605_));
 OAI21_X1 _3048_ (.A(\coll_reg[1] ),
    .B1(\coll_reg[2] ),
    .B2(\coll_reg[3] ),
    .ZN(_1616_));
 NAND2_X1 _3049_ (.A1(_1561_),
    .A2(_1616_),
    .ZN(_1627_));
 XNOR2_X1 _3050_ (.A(_1605_),
    .B(_1627_),
    .ZN(_1638_));
 XNOR2_X1 _3051_ (.A(\coll_reg[1] ),
    .B(_1638_),
    .ZN(_1649_));
 OR2_X1 _3052_ (.A1(\coll_reg[3] ),
    .A2(\coll_reg[2] ),
    .ZN(_1660_));
 OAI22_X1 _3053_ (.A1(\coll_reg[0] ),
    .A2(_1572_),
    .B1(_1660_),
    .B2(\coll_reg[1] ),
    .ZN(_1671_));
 XOR2_X1 _3054_ (.A(_1649_),
    .B(_1671_),
    .Z(_1682_));
 XNOR2_X1 _3055_ (.A(_1583_),
    .B(_1682_),
    .ZN(_1693_));
 XNOR2_X1 _3056_ (.A(_0012_),
    .B(_1693_),
    .ZN(_1704_));
 XOR2_X1 _3057_ (.A(_1539_),
    .B(_1704_),
    .Z(_1715_));
 XNOR2_X1 _3058_ (.A(_0015_),
    .B(_1715_),
    .ZN(_1726_));
 XNOR2_X1 _3059_ (.A(_1517_),
    .B(_1726_),
    .ZN(_1737_));
 XNOR2_X1 _3060_ (.A(_1506_),
    .B(_1737_),
    .ZN(_1748_));
 XNOR2_X1 _3061_ (.A(_1484_),
    .B(_1748_),
    .ZN(_1759_));
 XNOR2_X1 _3062_ (.A(\section_2.xn2[3] ),
    .B(_1759_),
    .ZN(_1770_));
 NAND2_X1 _3063_ (.A1(_1473_),
    .A2(_1770_),
    .ZN(_1781_));
 XNOR2_X1 _3064_ (.A(_1473_),
    .B(_1770_),
    .ZN(_1792_));
 XNOR2_X1 _3065_ (.A(\section_2.xn2[1] ),
    .B(\section_2.xn2[2] ),
    .ZN(_1803_));
 OAI21_X1 _3066_ (.A(_1781_),
    .B1(_1792_),
    .B2(_1803_),
    .ZN(_1814_));
 OAI22_X1 _3067_ (.A1(_0019_),
    .A2(_1748_),
    .B1(_1759_),
    .B2(_1440_),
    .ZN(_1825_));
 OR2_X1 _3068_ (.A1(_1539_),
    .A2(_1704_),
    .ZN(_1836_));
 NAND2_X1 _3069_ (.A1(_0015_),
    .A2(_1715_),
    .ZN(_1847_));
 NAND2_X1 _3070_ (.A1(_1836_),
    .A2(_1847_),
    .ZN(_1858_));
 NOR2_X1 _3071_ (.A1(\section_1.yn2[3] ),
    .A2(_1693_),
    .ZN(_1869_));
 NAND3_X1 _3072_ (.A1(\coll_reg[0] ),
    .A2(_1572_),
    .A3(_1649_),
    .ZN(_1880_));
 NOR2_X1 _3073_ (.A1(_1649_),
    .A2(_1671_),
    .ZN(_1891_));
 AOI21_X1 _3074_ (.A(_1605_),
    .B1(_1616_),
    .B2(_1561_),
    .ZN(_1902_));
 AOI21_X1 _3075_ (.A(_1902_),
    .B1(_1638_),
    .B2(\coll_reg[1] ),
    .ZN(_1913_));
 AND2_X1 _3076_ (.A1(\coll_reg[4] ),
    .A2(\coll_reg[3] ),
    .ZN(_1924_));
 AOI21_X1 _3077_ (.A(_1924_),
    .B1(_1594_),
    .B2(\coll_reg[2] ),
    .ZN(_1935_));
 XOR2_X1 _3078_ (.A(\coll_reg[5] ),
    .B(\coll_reg[3] ),
    .Z(_1946_));
 XNOR2_X1 _3079_ (.A(\coll_reg[4] ),
    .B(_1946_),
    .ZN(_1957_));
 XOR2_X1 _3080_ (.A(_1935_),
    .B(_1957_),
    .Z(_1968_));
 XNOR2_X1 _3081_ (.A(_1352_),
    .B(_1968_),
    .ZN(_1979_));
 XOR2_X1 _3082_ (.A(_1913_),
    .B(_1979_),
    .Z(_1990_));
 XOR2_X1 _3083_ (.A(_1891_),
    .B(_1990_),
    .Z(_2001_));
 XNOR2_X1 _3084_ (.A(_1880_),
    .B(_2001_),
    .ZN(_2012_));
 XNOR2_X1 _3085_ (.A(_0011_),
    .B(_2012_),
    .ZN(_2023_));
 XNOR2_X1 _3086_ (.A(_1869_),
    .B(_2023_),
    .ZN(_2034_));
 XNOR2_X1 _3087_ (.A(_0014_),
    .B(_2034_),
    .ZN(_2045_));
 XNOR2_X1 _3088_ (.A(_1858_),
    .B(_2045_),
    .ZN(_2056_));
 OR2_X1 _3089_ (.A1(_1517_),
    .A2(_1726_),
    .ZN(_2067_));
 OAI21_X1 _3090_ (.A(_2067_),
    .B1(_1737_),
    .B2(_1506_),
    .ZN(_2078_));
 XNOR2_X1 _3091_ (.A(_2056_),
    .B(_2078_),
    .ZN(_2089_));
 XOR2_X1 _3092_ (.A(\section_2.xn2[5] ),
    .B(_2089_),
    .Z(_2100_));
 XNOR2_X1 _3093_ (.A(\section_2.xn2[4] ),
    .B(_2100_),
    .ZN(_2111_));
 XNOR2_X1 _3094_ (.A(_1825_),
    .B(_2111_),
    .ZN(_2122_));
 XNOR2_X1 _3095_ (.A(\section_2.xn2[2] ),
    .B(\section_2.xn2[3] ),
    .ZN(_2133_));
 XOR2_X1 _3096_ (.A(_2122_),
    .B(_2133_),
    .Z(_2144_));
 NAND2_X1 _3097_ (.A1(_1814_),
    .A2(_2144_),
    .ZN(_2155_));
 XNOR2_X1 _3098_ (.A(_1814_),
    .B(_2144_),
    .ZN(_2166_));
 NAND2_X1 _3099_ (.A1(\section_2.xn2[1] ),
    .A2(\section_2.xn2[2] ),
    .ZN(_2177_));
 XNOR2_X1 _3100_ (.A(_0024_),
    .B(_2177_),
    .ZN(_2188_));
 OAI21_X1 _3101_ (.A(_2155_),
    .B1(_2166_),
    .B2(_2188_),
    .ZN(_2199_));
 NAND2_X1 _3102_ (.A1(_1825_),
    .A2(_2111_),
    .ZN(_2210_));
 OAI21_X1 _3103_ (.A(_2210_),
    .B1(_2122_),
    .B2(_2133_),
    .ZN(_2221_));
 OAI22_X1 _3104_ (.A1(_0017_),
    .A2(_2089_),
    .B1(_2100_),
    .B2(_1484_),
    .ZN(_2232_));
 INV_X1 _3105_ (.A(\section_2.xn2[6] ),
    .ZN(_2240_));
 OAI21_X1 _3106_ (.A(_2023_),
    .B1(_1693_),
    .B2(\section_1.yn2[3] ),
    .ZN(_2246_));
 NAND2_X1 _3107_ (.A1(_0014_),
    .A2(_2034_),
    .ZN(_2256_));
 NAND2_X1 _3108_ (.A1(_2246_),
    .A2(_2256_),
    .ZN(_2267_));
 NAND2_X1 _3109_ (.A1(\section_1.yn2[4] ),
    .A2(_2012_),
    .ZN(_2274_));
 INV_X1 _3110_ (.A(net86),
    .ZN(_2275_));
 NAND4_X1 _3111_ (.A1(\coll_reg[0] ),
    .A2(_1572_),
    .A3(_1649_),
    .A4(_1990_),
    .ZN(_2276_));
 AND2_X1 _3112_ (.A1(\coll_reg[2] ),
    .A2(\coll_reg[0] ),
    .ZN(_2277_));
 NOR2_X1 _3113_ (.A1(_1935_),
    .A2(_1957_),
    .ZN(_2278_));
 AOI21_X1 _3114_ (.A(_2278_),
    .B1(_1968_),
    .B2(_1352_),
    .ZN(_2279_));
 XOR2_X1 _3115_ (.A(\coll_reg[3] ),
    .B(\coll_reg[1] ),
    .Z(_2280_));
 NOR2_X1 _3116_ (.A1(\coll_reg[4] ),
    .A2(\coll_reg[3] ),
    .ZN(_2281_));
 NAND2_X1 _3117_ (.A1(\coll_reg[4] ),
    .A2(\coll_reg[3] ),
    .ZN(_2282_));
 INV_X1 _3118_ (.A(net87),
    .ZN(_2283_));
 AOI21_X1 _3119_ (.A(_2281_),
    .B1(_2282_),
    .B2(_2283_),
    .ZN(_2284_));
 XOR2_X1 _3120_ (.A(\coll_reg[6] ),
    .B(\coll_reg[5] ),
    .Z(_2285_));
 XNOR2_X1 _3121_ (.A(\coll_reg[4] ),
    .B(_2285_),
    .ZN(_2286_));
 XNOR2_X1 _3122_ (.A(_2284_),
    .B(_2286_),
    .ZN(_2287_));
 XNOR2_X1 _3123_ (.A(_2280_),
    .B(_2287_),
    .ZN(_2288_));
 XOR2_X1 _3124_ (.A(_2279_),
    .B(_2288_),
    .Z(_2289_));
 XOR2_X1 _3125_ (.A(_2277_),
    .B(_2289_),
    .Z(_2290_));
 NOR2_X1 _3126_ (.A1(_1913_),
    .A2(_1979_),
    .ZN(_2291_));
 AOI21_X1 _3127_ (.A(_2291_),
    .B1(_1990_),
    .B2(_1891_),
    .ZN(_2292_));
 XOR2_X1 _3128_ (.A(_2290_),
    .B(_2292_),
    .Z(_2293_));
 XNOR2_X1 _3129_ (.A(_2276_),
    .B(_2293_),
    .ZN(_2294_));
 XNOR2_X1 _3130_ (.A(_2275_),
    .B(_2294_),
    .ZN(_2295_));
 XOR2_X1 _3131_ (.A(_2274_),
    .B(_2295_),
    .Z(_2296_));
 XNOR2_X1 _3132_ (.A(\section_1.yn2[2] ),
    .B(_2296_),
    .ZN(_2297_));
 XOR2_X1 _3133_ (.A(_2267_),
    .B(_2297_),
    .Z(_2298_));
 AOI21_X1 _3134_ (.A(_2045_),
    .B1(_1847_),
    .B2(_1836_),
    .ZN(_2299_));
 AOI21_X1 _3135_ (.A(_2299_),
    .B1(_2056_),
    .B2(_2078_),
    .ZN(_2300_));
 XNOR2_X1 _3136_ (.A(_2298_),
    .B(_2300_),
    .ZN(_2301_));
 XNOR2_X1 _3137_ (.A(_2240_),
    .B(_2301_),
    .ZN(_2302_));
 XOR2_X1 _3138_ (.A(\section_2.xn2[5] ),
    .B(_2302_),
    .Z(_2303_));
 XNOR2_X1 _3139_ (.A(_2232_),
    .B(_2303_),
    .ZN(_2304_));
 XNOR2_X1 _3140_ (.A(\section_2.xn2[3] ),
    .B(\section_2.xn2[4] ),
    .ZN(_2305_));
 XOR2_X1 _3141_ (.A(_2304_),
    .B(_2305_),
    .Z(_2306_));
 XNOR2_X1 _3142_ (.A(_2221_),
    .B(_2306_),
    .ZN(_2307_));
 NAND2_X1 _3143_ (.A1(\section_2.xn2[2] ),
    .A2(\section_2.xn2[3] ),
    .ZN(_2308_));
 XOR2_X1 _3144_ (.A(_0023_),
    .B(_2308_),
    .Z(_2309_));
 XNOR2_X1 _3145_ (.A(_2307_),
    .B(_2309_),
    .ZN(_2310_));
 NAND2_X1 _3146_ (.A1(_2199_),
    .A2(_2310_),
    .ZN(_2311_));
 XNOR2_X1 _3147_ (.A(_2199_),
    .B(_2310_),
    .ZN(_2312_));
 OR2_X1 _3148_ (.A1(_0024_),
    .A2(_2177_),
    .ZN(_2313_));
 OAI21_X1 _3149_ (.A(_2311_),
    .B1(_2312_),
    .B2(_2313_),
    .ZN(_2314_));
 OR2_X1 _3150_ (.A1(_0023_),
    .A2(_2308_),
    .ZN(_2315_));
 NAND2_X1 _3151_ (.A1(_2221_),
    .A2(_2306_),
    .ZN(_2316_));
 INV_X1 _3152_ (.A(_2309_),
    .ZN(_2317_));
 OAI21_X1 _3153_ (.A(_2316_),
    .B1(_2307_),
    .B2(_2317_),
    .ZN(_2318_));
 NAND2_X1 _3154_ (.A1(_2232_),
    .A2(_2303_),
    .ZN(_2319_));
 OAI21_X1 _3155_ (.A(_2319_),
    .B1(_2304_),
    .B2(_2305_),
    .ZN(_2320_));
 AND2_X1 _3156_ (.A1(\section_2.xn2[5] ),
    .A2(_2302_),
    .ZN(_2321_));
 INV_X1 _3157_ (.A(_0020_),
    .ZN(_2322_));
 AND2_X1 _3158_ (.A1(_2322_),
    .A2(_2301_),
    .ZN(_2323_));
 NOR2_X1 _3159_ (.A1(_2321_),
    .A2(_2323_),
    .ZN(_2324_));
 INV_X1 _3160_ (.A(\section_2.xn2[7] ),
    .ZN(_2325_));
 NAND2_X1 _3161_ (.A1(_2267_),
    .A2(_2297_),
    .ZN(_2326_));
 NOR2_X1 _3162_ (.A1(_2275_),
    .A2(_2294_),
    .ZN(_2327_));
 INV_X1 _3163_ (.A(net63),
    .ZN(_2328_));
 NAND3_X1 _3164_ (.A1(_1891_),
    .A2(_1990_),
    .A3(_2290_),
    .ZN(_2329_));
 OAI21_X1 _3165_ (.A(_2329_),
    .B1(_2293_),
    .B2(_2276_),
    .ZN(_2330_));
 NAND2_X1 _3166_ (.A1(_2291_),
    .A2(_2290_),
    .ZN(_2331_));
 NOR2_X1 _3167_ (.A1(_2279_),
    .A2(_2288_),
    .ZN(_2332_));
 AOI21_X1 _3168_ (.A(_2332_),
    .B1(_2289_),
    .B2(_2277_),
    .ZN(_2333_));
 NAND2_X1 _3169_ (.A1(\coll_reg[3] ),
    .A2(\coll_reg[1] ),
    .ZN(_2334_));
 INV_X1 _3170_ (.A(_2334_),
    .ZN(_2335_));
 AOI211_X1 _3171_ (.A(_2281_),
    .B(_2286_),
    .C1(_2282_),
    .C2(_2283_),
    .ZN(_2336_));
 AOI21_X1 _3172_ (.A(_2336_),
    .B1(_2287_),
    .B2(_2280_),
    .ZN(_2337_));
 AND2_X1 _3173_ (.A1(\coll_reg[6] ),
    .A2(\coll_reg[5] ),
    .ZN(_2338_));
 AOI21_X1 _3174_ (.A(_2338_),
    .B1(_2285_),
    .B2(\coll_reg[4] ),
    .ZN(_2339_));
 XOR2_X1 _3175_ (.A(\coll_reg[7] ),
    .B(\coll_reg[6] ),
    .Z(_2340_));
 XNOR2_X1 _3176_ (.A(_0007_),
    .B(_2340_),
    .ZN(_2341_));
 XOR2_X1 _3177_ (.A(_2339_),
    .B(_2341_),
    .Z(_2342_));
 OR2_X1 _3178_ (.A1(\coll_reg[4] ),
    .A2(\coll_reg[2] ),
    .ZN(_2343_));
 NAND2_X1 _3179_ (.A1(\coll_reg[4] ),
    .A2(\coll_reg[2] ),
    .ZN(_2344_));
 NAND2_X1 _3180_ (.A1(_2343_),
    .A2(_2344_),
    .ZN(_2345_));
 XNOR2_X1 _3181_ (.A(_2342_),
    .B(_2345_),
    .ZN(_2346_));
 XOR2_X1 _3182_ (.A(_2337_),
    .B(_2346_),
    .Z(_2347_));
 XNOR2_X1 _3183_ (.A(_2335_),
    .B(_2347_),
    .ZN(_2348_));
 XNOR2_X1 _3184_ (.A(_2333_),
    .B(_2348_),
    .ZN(_2349_));
 XOR2_X1 _3185_ (.A(_2331_),
    .B(_2349_),
    .Z(_2350_));
 XOR2_X1 _3186_ (.A(_2330_),
    .B(_2350_),
    .Z(_2351_));
 XNOR2_X1 _3187_ (.A(_2328_),
    .B(_2351_),
    .ZN(_2352_));
 XOR2_X1 _3188_ (.A(_2327_),
    .B(_2352_),
    .Z(_2353_));
 XNOR2_X1 _3189_ (.A(\section_1.yn2[3] ),
    .B(_2353_),
    .ZN(_2354_));
 NOR2_X1 _3190_ (.A1(_2274_),
    .A2(_2295_),
    .ZN(_2355_));
 AOI21_X1 _3191_ (.A(_2355_),
    .B1(_2296_),
    .B2(_0013_),
    .ZN(_2356_));
 XOR2_X1 _3192_ (.A(_2354_),
    .B(_2356_),
    .Z(_2357_));
 XOR2_X1 _3193_ (.A(_2326_),
    .B(_2357_),
    .Z(_2358_));
 INV_X1 _3194_ (.A(_2298_),
    .ZN(_2359_));
 NOR2_X1 _3195_ (.A1(_2359_),
    .A2(_2300_),
    .ZN(_2360_));
 XNOR2_X1 _3196_ (.A(_2358_),
    .B(_2360_),
    .ZN(_2361_));
 XNOR2_X1 _3197_ (.A(_2325_),
    .B(_2361_),
    .ZN(_2362_));
 XNOR2_X1 _3198_ (.A(\section_2.xn2[6] ),
    .B(_2362_),
    .ZN(_2363_));
 XNOR2_X1 _3199_ (.A(_2324_),
    .B(_2363_),
    .ZN(_2364_));
 XOR2_X1 _3200_ (.A(\section_2.xn2[4] ),
    .B(\section_2.xn2[5] ),
    .Z(_2365_));
 XNOR2_X1 _3201_ (.A(_2364_),
    .B(_2365_),
    .ZN(_2366_));
 XOR2_X1 _3202_ (.A(_2320_),
    .B(_2366_),
    .Z(_2367_));
 NAND2_X1 _3203_ (.A1(\section_2.xn2[3] ),
    .A2(\section_2.xn2[4] ),
    .ZN(_2368_));
 XOR2_X1 _3204_ (.A(_0022_),
    .B(_2368_),
    .Z(_2369_));
 XNOR2_X1 _3205_ (.A(_2367_),
    .B(_2369_),
    .ZN(_2370_));
 XNOR2_X1 _3206_ (.A(_2318_),
    .B(_2370_),
    .ZN(_2371_));
 XOR2_X1 _3207_ (.A(_2315_),
    .B(_2371_),
    .Z(_2372_));
 AND2_X1 _3208_ (.A1(_2314_),
    .A2(_2372_),
    .ZN(_2373_));
 XOR2_X1 _3209_ (.A(_2314_),
    .B(_2372_),
    .Z(_2374_));
 XNOR2_X1 _3210_ (.A(\section_2.xn2[0] ),
    .B(\section_2.xn2[1] ),
    .ZN(_2375_));
 XNOR2_X1 _3211_ (.A(_1462_),
    .B(_1451_),
    .ZN(_2376_));
 XNOR2_X1 _3212_ (.A(_1396_),
    .B(_1407_),
    .ZN(_2377_));
 OR2_X1 _3213_ (.A1(_0022_),
    .A2(_2377_),
    .ZN(_2378_));
 XNOR2_X1 _3214_ (.A(_1462_),
    .B(_2377_),
    .ZN(_2379_));
 INV_X1 _3215_ (.A(_2379_),
    .ZN(_2380_));
 NAND2_X1 _3216_ (.A1(\section_2.xn2[1] ),
    .A2(_2380_),
    .ZN(_2381_));
 AOI21_X1 _3217_ (.A(_2376_),
    .B1(_2378_),
    .B2(_2381_),
    .ZN(_2382_));
 AND3_X1 _3218_ (.A1(_2381_),
    .A2(_2378_),
    .A3(_2376_),
    .ZN(_2383_));
 OR2_X1 _3219_ (.A1(_2382_),
    .A2(_2383_),
    .ZN(_2384_));
 XNOR2_X1 _3220_ (.A(_2375_),
    .B(_2384_),
    .ZN(_2385_));
 INV_X1 _3221_ (.A(net41),
    .ZN(_2386_));
 XNOR2_X1 _3222_ (.A(_2386_),
    .B(_1385_),
    .ZN(_2387_));
 INV_X1 _3223_ (.A(_2387_),
    .ZN(_2388_));
 XNOR2_X1 _3224_ (.A(\section_2.xn2[1] ),
    .B(_2387_),
    .ZN(_2389_));
 INV_X1 _3225_ (.A(\section_2.xn2[0] ),
    .ZN(_2390_));
 OAI22_X1 _3226_ (.A1(_0023_),
    .A2(_2388_),
    .B1(_2389_),
    .B2(_2390_),
    .ZN(_2391_));
 XNOR2_X1 _3227_ (.A(\section_2.xn2[1] ),
    .B(_2379_),
    .ZN(_2392_));
 AND2_X1 _3228_ (.A1(_2391_),
    .A2(_2392_),
    .ZN(_2393_));
 XOR2_X1 _3229_ (.A(_2391_),
    .B(_2392_),
    .Z(_2394_));
 AOI21_X1 _3230_ (.A(_2393_),
    .B1(_2394_),
    .B2(\section_2.xn2[0] ),
    .ZN(_2395_));
 NOR2_X1 _3231_ (.A1(_2385_),
    .A2(_2395_),
    .ZN(_2396_));
 NAND2_X1 _3232_ (.A1(\section_2.xn2[0] ),
    .A2(\section_2.xn2[1] ),
    .ZN(_2397_));
 NOR2_X1 _3233_ (.A1(_2375_),
    .A2(_2384_),
    .ZN(_2398_));
 NOR2_X1 _3234_ (.A1(_2382_),
    .A2(_2398_),
    .ZN(_2399_));
 XOR2_X1 _3235_ (.A(_1792_),
    .B(_1803_),
    .Z(_2400_));
 XNOR2_X1 _3236_ (.A(_2399_),
    .B(_2400_),
    .ZN(_2401_));
 XNOR2_X1 _3237_ (.A(_2397_),
    .B(_2401_),
    .ZN(_2402_));
 OAI21_X1 _3238_ (.A(_2400_),
    .B1(_2398_),
    .B2(_2382_),
    .ZN(_2403_));
 NAND3_X1 _3239_ (.A1(\section_2.xn2[0] ),
    .A2(\section_2.xn2[1] ),
    .A3(_2401_),
    .ZN(_2404_));
 NAND2_X1 _3240_ (.A1(_2403_),
    .A2(_2404_),
    .ZN(_2405_));
 XOR2_X1 _3241_ (.A(_2166_),
    .B(_2188_),
    .Z(_2406_));
 XOR2_X1 _3242_ (.A(_2405_),
    .B(_2406_),
    .Z(_2407_));
 NAND3_X1 _3243_ (.A1(_2396_),
    .A2(_2402_),
    .A3(_2407_),
    .ZN(_2408_));
 NAND3_X1 _3244_ (.A1(\coll_reg[0] ),
    .A2(\section_2.xn2[0] ),
    .A3(_2389_),
    .ZN(_2409_));
 NOR2_X1 _3245_ (.A1(_2394_),
    .A2(_2409_),
    .ZN(_2410_));
 XOR2_X1 _3246_ (.A(_2385_),
    .B(_2395_),
    .Z(_2411_));
 NAND2_X1 _3247_ (.A1(_2410_),
    .A2(_2411_),
    .ZN(_2412_));
 XNOR2_X1 _3248_ (.A(_2396_),
    .B(_2402_),
    .ZN(_2413_));
 OR2_X1 _3249_ (.A1(_2412_),
    .A2(_2413_),
    .ZN(_2414_));
 NAND2_X1 _3250_ (.A1(_2396_),
    .A2(_2402_),
    .ZN(_2415_));
 XNOR2_X1 _3251_ (.A(_2415_),
    .B(_2407_),
    .ZN(_2416_));
 INV_X1 _3252_ (.A(_2416_),
    .ZN(_2417_));
 OAI21_X1 _3253_ (.A(_2408_),
    .B1(_2414_),
    .B2(_2417_),
    .ZN(_2418_));
 NAND2_X1 _3254_ (.A1(_2405_),
    .A2(_2406_),
    .ZN(_2419_));
 XOR2_X1 _3255_ (.A(_2313_),
    .B(_2312_),
    .Z(_2420_));
 XNOR2_X1 _3256_ (.A(_2419_),
    .B(_2420_),
    .ZN(_2421_));
 NAND2_X1 _3257_ (.A1(_2418_),
    .A2(_2421_),
    .ZN(_2422_));
 INV_X1 _3258_ (.A(_2420_),
    .ZN(_2423_));
 OAI21_X1 _3259_ (.A(_2422_),
    .B1(_2423_),
    .B2(_2419_),
    .ZN(_2424_));
 AOI21_X1 _3260_ (.A(_2373_),
    .B1(_2374_),
    .B2(_2424_),
    .ZN(_2425_));
 NAND2_X1 _3261_ (.A1(_2318_),
    .A2(_2370_),
    .ZN(_2426_));
 OAI21_X1 _3262_ (.A(_2426_),
    .B1(_2371_),
    .B2(_2315_),
    .ZN(_2427_));
 NOR2_X1 _3263_ (.A1(_0022_),
    .A2(_2368_),
    .ZN(_2428_));
 INV_X1 _3264_ (.A(_2366_),
    .ZN(_2429_));
 NAND2_X1 _3265_ (.A1(_2320_),
    .A2(_2429_),
    .ZN(_2430_));
 INV_X1 _3266_ (.A(_2369_),
    .ZN(_2431_));
 OR2_X1 _3267_ (.A1(_2367_),
    .A2(_2431_),
    .ZN(_2432_));
 NAND2_X1 _3268_ (.A1(_2430_),
    .A2(_2432_),
    .ZN(_2433_));
 OAI21_X1 _3269_ (.A(_2363_),
    .B1(_2323_),
    .B2(_2321_),
    .ZN(_2434_));
 NAND2_X1 _3270_ (.A1(_2364_),
    .A2(_2365_),
    .ZN(_2435_));
 NAND2_X1 _3271_ (.A1(_2434_),
    .A2(_2435_),
    .ZN(_2436_));
 OAI22_X1 _3272_ (.A1(_0018_),
    .A2(_2361_),
    .B1(_2362_),
    .B2(_2240_),
    .ZN(_2437_));
 NOR2_X1 _3273_ (.A1(_2326_),
    .A2(_2357_),
    .ZN(_2438_));
 AOI21_X1 _3274_ (.A(_2438_),
    .B1(_2358_),
    .B2(_2360_),
    .ZN(_2439_));
 INV_X1 _3275_ (.A(_2354_),
    .ZN(_2440_));
 NOR2_X1 _3276_ (.A1(_2440_),
    .A2(_2356_),
    .ZN(_2441_));
 NAND2_X1 _3277_ (.A1(\section_1.yn2[6] ),
    .A2(_2351_),
    .ZN(_2442_));
 INV_X1 _3278_ (.A(net85),
    .ZN(_2443_));
 NOR2_X1 _3279_ (.A1(_2333_),
    .A2(_2348_),
    .ZN(_2444_));
 NOR2_X1 _3280_ (.A1(_2337_),
    .A2(_2346_),
    .ZN(_2445_));
 AOI21_X1 _3281_ (.A(_2445_),
    .B1(_2347_),
    .B2(_2335_),
    .ZN(_2446_));
 AND2_X1 _3282_ (.A1(\coll_reg[4] ),
    .A2(_2285_),
    .ZN(_2447_));
 OAI21_X1 _3283_ (.A(_2341_),
    .B1(_2447_),
    .B2(_2338_),
    .ZN(_2448_));
 OAI21_X1 _3284_ (.A(_2448_),
    .B1(_2342_),
    .B2(_2345_),
    .ZN(_2449_));
 XOR2_X1 _3285_ (.A(\coll_reg[8] ),
    .B(\coll_reg[7] ),
    .Z(_2450_));
 XNOR2_X1 _3286_ (.A(\coll_reg[6] ),
    .B(_2450_),
    .ZN(_2451_));
 NAND2_X1 _3287_ (.A1(\coll_reg[7] ),
    .A2(\coll_reg[6] ),
    .ZN(_2452_));
 OAI21_X1 _3288_ (.A(\coll_reg[5] ),
    .B1(\coll_reg[6] ),
    .B2(\coll_reg[7] ),
    .ZN(_2453_));
 NAND2_X1 _3289_ (.A1(_2452_),
    .A2(_2453_),
    .ZN(_2454_));
 XNOR2_X1 _3290_ (.A(_2451_),
    .B(_2454_),
    .ZN(_2455_));
 XOR2_X1 _3291_ (.A(_1946_),
    .B(_2455_),
    .Z(_2456_));
 XNOR2_X1 _3292_ (.A(_2449_),
    .B(_2456_),
    .ZN(_2457_));
 XNOR2_X1 _3293_ (.A(_2344_),
    .B(_2457_),
    .ZN(_2458_));
 XOR2_X1 _3294_ (.A(_2446_),
    .B(_2458_),
    .Z(_2459_));
 NAND2_X1 _3295_ (.A1(_2444_),
    .A2(_2459_),
    .ZN(_2460_));
 OR2_X1 _3296_ (.A1(_2444_),
    .A2(_2459_),
    .ZN(_2461_));
 NAND2_X1 _3297_ (.A1(_2460_),
    .A2(_2461_),
    .ZN(_2462_));
 NOR2_X1 _3298_ (.A1(_2331_),
    .A2(_2349_),
    .ZN(_2463_));
 AOI21_X1 _3299_ (.A(_2463_),
    .B1(_2350_),
    .B2(_2330_),
    .ZN(_2464_));
 XNOR2_X1 _3300_ (.A(_2462_),
    .B(_2464_),
    .ZN(_2465_));
 XNOR2_X1 _3301_ (.A(_2443_),
    .B(_2465_),
    .ZN(_2466_));
 XOR2_X1 _3302_ (.A(_2442_),
    .B(_2466_),
    .Z(_2467_));
 XNOR2_X1 _3303_ (.A(\section_1.yn2[4] ),
    .B(_2467_),
    .ZN(_2468_));
 AND2_X1 _3304_ (.A1(_2327_),
    .A2(_2352_),
    .ZN(_2469_));
 AOI21_X1 _3305_ (.A(_2469_),
    .B1(_2353_),
    .B2(_0012_),
    .ZN(_2470_));
 XNOR2_X1 _3306_ (.A(_2468_),
    .B(_2470_),
    .ZN(_2471_));
 XNOR2_X1 _3307_ (.A(_2441_),
    .B(_2471_),
    .ZN(_2472_));
 XOR2_X1 _3308_ (.A(_2439_),
    .B(_2472_),
    .Z(_2473_));
 XNOR2_X1 _3309_ (.A(\section_2.xn2[8] ),
    .B(_2473_),
    .ZN(_2474_));
 XOR2_X1 _3310_ (.A(_0018_),
    .B(_2474_),
    .Z(_2475_));
 XNOR2_X1 _3311_ (.A(_2437_),
    .B(_2475_),
    .ZN(_2476_));
 XNOR2_X1 _3312_ (.A(\section_2.xn2[5] ),
    .B(\section_2.xn2[6] ),
    .ZN(_2477_));
 XNOR2_X1 _3313_ (.A(_2476_),
    .B(_2477_),
    .ZN(_2478_));
 XNOR2_X1 _3314_ (.A(_2436_),
    .B(_2478_),
    .ZN(_2479_));
 NAND2_X1 _3315_ (.A1(\section_2.xn2[4] ),
    .A2(\section_2.xn2[5] ),
    .ZN(_2480_));
 XOR2_X1 _3316_ (.A(_0021_),
    .B(_2480_),
    .Z(_2481_));
 XNOR2_X1 _3317_ (.A(_2479_),
    .B(_2481_),
    .ZN(_2482_));
 XOR2_X1 _3318_ (.A(_2433_),
    .B(_2482_),
    .Z(_2483_));
 XNOR2_X1 _3319_ (.A(_2428_),
    .B(_2483_),
    .ZN(_2484_));
 XNOR2_X1 _3320_ (.A(_2427_),
    .B(_2484_),
    .ZN(_2485_));
 XOR2_X1 _3321_ (.A(_2425_),
    .B(_2485_),
    .Z(_2486_));
 NAND2_X1 _3322_ (.A1(z[5]),
    .A2(_2486_),
    .ZN(_2487_));
 AOI21_X1 _3323_ (.A(_2482_),
    .B1(_2432_),
    .B2(_2430_),
    .ZN(_2488_));
 NAND3_X1 _3324_ (.A1(_2430_),
    .A2(_2432_),
    .A3(_2482_),
    .ZN(_2489_));
 AOI21_X1 _3325_ (.A(_2488_),
    .B1(_2489_),
    .B2(_2428_),
    .ZN(_2490_));
 NOR2_X1 _3326_ (.A1(_0021_),
    .A2(_2480_),
    .ZN(_2491_));
 AOI21_X1 _3327_ (.A(_2478_),
    .B1(_2435_),
    .B2(_2434_),
    .ZN(_2492_));
 AOI21_X1 _3328_ (.A(_2492_),
    .B1(_2479_),
    .B2(_2481_),
    .ZN(_2493_));
 NAND2_X1 _3329_ (.A1(_2437_),
    .A2(_2475_),
    .ZN(_2494_));
 NOR2_X1 _3330_ (.A1(_2437_),
    .A2(_2475_),
    .ZN(_2495_));
 OAI21_X1 _3331_ (.A(_2494_),
    .B1(_2477_),
    .B2(_2495_),
    .ZN(_2496_));
 INV_X1 _3332_ (.A(_2473_),
    .ZN(_2497_));
 OAI22_X1 _3333_ (.A1(_0016_),
    .A2(_2497_),
    .B1(_2474_),
    .B2(_2325_),
    .ZN(_2498_));
 NAND2_X1 _3334_ (.A1(_2441_),
    .A2(_2471_),
    .ZN(_2499_));
 OAI21_X1 _3335_ (.A(_2499_),
    .B1(_2472_),
    .B2(_2439_),
    .ZN(_2500_));
 INV_X1 _3336_ (.A(_2470_),
    .ZN(_2501_));
 NAND2_X1 _3337_ (.A1(_2468_),
    .A2(_2501_),
    .ZN(_2502_));
 OR2_X1 _3338_ (.A1(_2443_),
    .A2(_2465_),
    .ZN(_2503_));
 INV_X1 _3339_ (.A(net77),
    .ZN(_2504_));
 NOR2_X1 _3340_ (.A1(_2446_),
    .A2(_2458_),
    .ZN(_2505_));
 NAND2_X1 _3341_ (.A1(_2449_),
    .A2(_2456_),
    .ZN(_2506_));
 OAI21_X1 _3342_ (.A(_2506_),
    .B1(_2457_),
    .B2(_2344_),
    .ZN(_2507_));
 NOR2_X1 _3343_ (.A1(_2283_),
    .A2(_1286_),
    .ZN(_2508_));
 AOI21_X1 _3344_ (.A(_2451_),
    .B1(_2453_),
    .B2(_2452_),
    .ZN(_2509_));
 AOI21_X1 _3345_ (.A(_2509_),
    .B1(_2455_),
    .B2(_1946_),
    .ZN(_2510_));
 AND2_X1 _3346_ (.A1(\coll_reg[8] ),
    .A2(\coll_reg[7] ),
    .ZN(_2511_));
 AOI21_X1 _3347_ (.A(_2511_),
    .B1(_2450_),
    .B2(\coll_reg[6] ),
    .ZN(_2512_));
 XOR2_X1 _3348_ (.A(\coll_reg[9] ),
    .B(\coll_reg[8] ),
    .Z(_2513_));
 XNOR2_X1 _3349_ (.A(\coll_reg[7] ),
    .B(_2513_),
    .ZN(_2514_));
 XOR2_X1 _3350_ (.A(_2512_),
    .B(_2514_),
    .Z(_2515_));
 XNOR2_X1 _3351_ (.A(\coll_reg[6] ),
    .B(\coll_reg[4] ),
    .ZN(_2516_));
 INV_X1 _3352_ (.A(_2516_),
    .ZN(_2517_));
 XNOR2_X1 _3353_ (.A(_2515_),
    .B(_2517_),
    .ZN(_2518_));
 XOR2_X1 _3354_ (.A(_2510_),
    .B(_2518_),
    .Z(_2519_));
 XOR2_X1 _3355_ (.A(_2508_),
    .B(_2519_),
    .Z(_2520_));
 XNOR2_X1 _3356_ (.A(_2507_),
    .B(_2520_),
    .ZN(_2521_));
 XNOR2_X1 _3357_ (.A(_2505_),
    .B(_2521_),
    .ZN(_2522_));
 OAI21_X1 _3358_ (.A(_2460_),
    .B1(_2462_),
    .B2(_2464_),
    .ZN(_2523_));
 XNOR2_X1 _3359_ (.A(_2522_),
    .B(_2523_),
    .ZN(_2524_));
 XNOR2_X1 _3360_ (.A(_2504_),
    .B(_2524_),
    .ZN(_2525_));
 XOR2_X1 _3361_ (.A(_2503_),
    .B(_2525_),
    .Z(_2526_));
 XNOR2_X1 _3362_ (.A(_0009_),
    .B(_2526_),
    .ZN(_2527_));
 NOR2_X1 _3363_ (.A1(_2442_),
    .A2(_2466_),
    .ZN(_2528_));
 AOI21_X1 _3364_ (.A(_2528_),
    .B1(_2467_),
    .B2(_0011_),
    .ZN(_2529_));
 XNOR2_X1 _3365_ (.A(_2527_),
    .B(_2529_),
    .ZN(_2530_));
 XOR2_X1 _3366_ (.A(_2502_),
    .B(_2530_),
    .Z(_2531_));
 XNOR2_X1 _3367_ (.A(_2500_),
    .B(_2531_),
    .ZN(_2532_));
 XNOR2_X1 _3368_ (.A(_0016_),
    .B(\section_2.xn2[9] ),
    .ZN(_2533_));
 XNOR2_X1 _3369_ (.A(_2532_),
    .B(_2533_),
    .ZN(_2534_));
 XNOR2_X1 _3370_ (.A(_2498_),
    .B(_2534_),
    .ZN(_2535_));
 XNOR2_X1 _3371_ (.A(\section_2.xn2[7] ),
    .B(\section_2.xn2[6] ),
    .ZN(_2536_));
 XOR2_X1 _3372_ (.A(_2535_),
    .B(_2536_),
    .Z(_2537_));
 XNOR2_X1 _3373_ (.A(_2496_),
    .B(_2537_),
    .ZN(_2538_));
 NAND2_X1 _3374_ (.A1(\section_2.xn2[5] ),
    .A2(\section_2.xn2[6] ),
    .ZN(_2539_));
 XNOR2_X1 _3375_ (.A(_0019_),
    .B(_2539_),
    .ZN(_2540_));
 XOR2_X1 _3376_ (.A(_2538_),
    .B(_2540_),
    .Z(_2541_));
 XNOR2_X1 _3377_ (.A(_2493_),
    .B(_2541_),
    .ZN(_2542_));
 XNOR2_X1 _3378_ (.A(_2491_),
    .B(_2542_),
    .ZN(_2543_));
 XNOR2_X1 _3379_ (.A(_2490_),
    .B(_2543_),
    .ZN(_2544_));
 NAND2_X1 _3380_ (.A1(_2427_),
    .A2(_2484_),
    .ZN(_2545_));
 OAI21_X1 _3381_ (.A(_2545_),
    .B1(_2485_),
    .B2(_2425_),
    .ZN(_2546_));
 XNOR2_X1 _3382_ (.A(_2544_),
    .B(_2546_),
    .ZN(_2547_));
 XNOR2_X1 _3383_ (.A(z[6]),
    .B(_2547_),
    .ZN(_2548_));
 NOR2_X1 _3384_ (.A1(_2487_),
    .A2(_2548_),
    .ZN(_2549_));
 NAND2_X1 _3385_ (.A1(z[6]),
    .A2(_2547_),
    .ZN(_2550_));
 NOR3_X1 _3386_ (.A1(_2425_),
    .A2(_2485_),
    .A3(_2544_),
    .ZN(_2551_));
 OR2_X1 _3387_ (.A1(_2490_),
    .A2(_2543_),
    .ZN(_2552_));
 OAI21_X1 _3388_ (.A(_2552_),
    .B1(_2544_),
    .B2(_2545_),
    .ZN(_2553_));
 OR2_X1 _3389_ (.A1(_2551_),
    .A2(_2553_),
    .ZN(_2554_));
 INV_X1 _3390_ (.A(_2541_),
    .ZN(_2555_));
 NOR2_X1 _3391_ (.A1(_2493_),
    .A2(_2555_),
    .ZN(_2556_));
 AOI21_X1 _3392_ (.A(_2556_),
    .B1(_2542_),
    .B2(_2491_),
    .ZN(_2557_));
 NOR2_X1 _3393_ (.A1(_0019_),
    .A2(_2539_),
    .ZN(_2558_));
 NOR2_X1 _3394_ (.A1(_2538_),
    .A2(_2540_),
    .ZN(_2559_));
 AOI21_X1 _3395_ (.A(_2559_),
    .B1(_2537_),
    .B2(_2496_),
    .ZN(_2560_));
 NAND2_X1 _3396_ (.A1(\section_2.xn2[7] ),
    .A2(\section_2.xn2[6] ),
    .ZN(_2561_));
 XOR2_X1 _3397_ (.A(_0017_),
    .B(_2561_),
    .Z(_2562_));
 NOR2_X1 _3398_ (.A1(_2535_),
    .A2(_2536_),
    .ZN(_2563_));
 AOI21_X1 _3399_ (.A(_2563_),
    .B1(_2534_),
    .B2(_2498_),
    .ZN(_2564_));
 XOR2_X1 _3400_ (.A(\section_2.xn2[8] ),
    .B(\section_2.xn2[7] ),
    .Z(_2565_));
 NOR2_X1 _3401_ (.A1(_2502_),
    .A2(_2530_),
    .ZN(_2566_));
 AOI21_X1 _3402_ (.A(_2566_),
    .B1(_2531_),
    .B2(_2500_),
    .ZN(_2567_));
 NOR2_X1 _3403_ (.A1(_2527_),
    .A2(_2529_),
    .ZN(_2568_));
 NOR2_X1 _3404_ (.A1(_2503_),
    .A2(_2525_),
    .ZN(_2569_));
 AOI21_X1 _3405_ (.A(_2569_),
    .B1(_2526_),
    .B2(_0009_),
    .ZN(_2570_));
 NOR2_X1 _3406_ (.A1(_0008_),
    .A2(_2524_),
    .ZN(_2571_));
 INV_X1 _3407_ (.A(net83),
    .ZN(_2572_));
 NOR3_X1 _3408_ (.A1(_2446_),
    .A2(_2458_),
    .A3(_2521_),
    .ZN(_2573_));
 AND2_X1 _3409_ (.A1(_2444_),
    .A2(_2459_),
    .ZN(_2574_));
 AOI21_X1 _3410_ (.A(_2573_),
    .B1(_2522_),
    .B2(_2574_),
    .ZN(_2575_));
 NAND3_X1 _3411_ (.A1(_2460_),
    .A2(_2461_),
    .A3(_2522_),
    .ZN(_2576_));
 OAI21_X1 _3412_ (.A(_2575_),
    .B1(_2576_),
    .B2(_2464_),
    .ZN(_2577_));
 NAND2_X1 _3413_ (.A1(_2507_),
    .A2(_2520_),
    .ZN(_2578_));
 NOR2_X1 _3414_ (.A1(_2510_),
    .A2(_2518_),
    .ZN(_2579_));
 AOI21_X1 _3415_ (.A(_2579_),
    .B1(_2519_),
    .B2(_2508_),
    .ZN(_2580_));
 AND2_X1 _3416_ (.A1(\coll_reg[6] ),
    .A2(\coll_reg[4] ),
    .ZN(_2581_));
 NOR2_X1 _3417_ (.A1(_2512_),
    .A2(_2514_),
    .ZN(_2582_));
 AOI21_X1 _3418_ (.A(_2582_),
    .B1(_2515_),
    .B2(_2517_),
    .ZN(_2583_));
 XNOR2_X1 _3419_ (.A(\coll_reg[7] ),
    .B(\coll_reg[5] ),
    .ZN(_2584_));
 INV_X1 _3420_ (.A(net92),
    .ZN(_2585_));
 XNOR2_X1 _3421_ (.A(\coll_reg[9] ),
    .B(\coll_reg[10] ),
    .ZN(_2586_));
 XNOR2_X1 _3422_ (.A(_2585_),
    .B(_2586_),
    .ZN(_2587_));
 AND2_X1 _3423_ (.A1(\coll_reg[9] ),
    .A2(\coll_reg[8] ),
    .ZN(_2588_));
 AOI21_X1 _3424_ (.A(_2588_),
    .B1(_2513_),
    .B2(\coll_reg[7] ),
    .ZN(_2589_));
 XNOR2_X1 _3425_ (.A(_2587_),
    .B(_2589_),
    .ZN(_2590_));
 XNOR2_X1 _3426_ (.A(_2584_),
    .B(_2590_),
    .ZN(_2591_));
 XOR2_X1 _3427_ (.A(_2583_),
    .B(_2591_),
    .Z(_2592_));
 XOR2_X1 _3428_ (.A(_2581_),
    .B(_2592_),
    .Z(_2593_));
 XOR2_X1 _3429_ (.A(_2580_),
    .B(_2593_),
    .Z(_2594_));
 XOR2_X1 _3430_ (.A(_2578_),
    .B(_2594_),
    .Z(_2595_));
 XNOR2_X1 _3431_ (.A(_2577_),
    .B(_2595_),
    .ZN(_2596_));
 XNOR2_X1 _3432_ (.A(_2572_),
    .B(_2596_),
    .ZN(_2597_));
 XNOR2_X1 _3433_ (.A(_2571_),
    .B(_2597_),
    .ZN(_2598_));
 XNOR2_X1 _3434_ (.A(_0003_),
    .B(_2598_),
    .ZN(_2599_));
 XOR2_X1 _3435_ (.A(_2570_),
    .B(_2599_),
    .Z(_2600_));
 XOR2_X1 _3436_ (.A(_2568_),
    .B(_2600_),
    .Z(_2601_));
 XNOR2_X1 _3437_ (.A(_2567_),
    .B(_2601_),
    .ZN(_2602_));
 XOR2_X1 _3438_ (.A(\section_2.xn2[10] ),
    .B(_2602_),
    .Z(_2603_));
 XNOR2_X1 _3439_ (.A(\section_2.xn2[9] ),
    .B(_2603_),
    .ZN(_2604_));
 NOR2_X1 _3440_ (.A1(\section_2.xn2[9] ),
    .A2(\section_2.xn2[8] ),
    .ZN(_2605_));
 NOR2_X1 _3441_ (.A1(_2532_),
    .A2(_2605_),
    .ZN(_2606_));
 AOI21_X1 _3442_ (.A(_2606_),
    .B1(\section_2.xn2[8] ),
    .B2(\section_2.xn2[9] ),
    .ZN(_2607_));
 XOR2_X1 _3443_ (.A(_2604_),
    .B(_2607_),
    .Z(_2608_));
 XNOR2_X1 _3444_ (.A(_2565_),
    .B(_2608_),
    .ZN(_2609_));
 XOR2_X1 _3445_ (.A(_2564_),
    .B(_2609_),
    .Z(_2610_));
 XNOR2_X1 _3446_ (.A(_2562_),
    .B(_2610_),
    .ZN(_2611_));
 XOR2_X1 _3447_ (.A(_2560_),
    .B(_2611_),
    .Z(_2612_));
 XNOR2_X1 _3448_ (.A(_2558_),
    .B(_2612_),
    .ZN(_2613_));
 XOR2_X1 _3449_ (.A(_2557_),
    .B(_2613_),
    .Z(_2614_));
 XOR2_X1 _3450_ (.A(_2554_),
    .B(_2614_),
    .Z(_2615_));
 XNOR2_X1 _3451_ (.A(z[7]),
    .B(_2615_),
    .ZN(_2616_));
 XOR2_X1 _3452_ (.A(_2550_),
    .B(_2616_),
    .Z(_2617_));
 XNOR2_X1 _3453_ (.A(_2549_),
    .B(_2617_),
    .ZN(_2618_));
 NOR2_X1 _3454_ (.A1(_1275_),
    .A2(_2618_),
    .ZN(_2619_));
 AOI21_X1 _3455_ (.A(_2619_),
    .B1(_2617_),
    .B2(_2549_),
    .ZN(_2620_));
 NAND2_X1 _3456_ (.A1(z[1]),
    .A2(z[0]),
    .ZN(_2621_));
 XOR2_X1 _3457_ (.A(z[2]),
    .B(z[1]),
    .Z(_2622_));
 XNOR2_X1 _3458_ (.A(_2621_),
    .B(_2622_),
    .ZN(_2623_));
 NOR2_X1 _3459_ (.A1(_2550_),
    .A2(_2616_),
    .ZN(_2624_));
 AND2_X1 _3460_ (.A1(z[7]),
    .A2(_2615_),
    .ZN(_2625_));
 INV_X1 _3461_ (.A(net79),
    .ZN(_2626_));
 NOR2_X1 _3462_ (.A1(_2557_),
    .A2(_2613_),
    .ZN(_2627_));
 AOI21_X1 _3463_ (.A(_2627_),
    .B1(_2614_),
    .B2(_2554_),
    .ZN(_2628_));
 NOR2_X1 _3464_ (.A1(_2560_),
    .A2(_2611_),
    .ZN(_2629_));
 AOI21_X1 _3465_ (.A(_2629_),
    .B1(_2612_),
    .B2(_2558_),
    .ZN(_2630_));
 NOR2_X1 _3466_ (.A1(_0017_),
    .A2(_2561_),
    .ZN(_2631_));
 NOR2_X1 _3467_ (.A1(_2564_),
    .A2(_2609_),
    .ZN(_2632_));
 AOI21_X1 _3468_ (.A(_2632_),
    .B1(_2610_),
    .B2(_2562_),
    .ZN(_2633_));
 NAND2_X1 _3469_ (.A1(\section_2.xn2[8] ),
    .A2(\section_2.xn2[7] ),
    .ZN(_2634_));
 XNOR2_X1 _3470_ (.A(_2322_),
    .B(_2634_),
    .ZN(_2635_));
 NOR2_X1 _3471_ (.A1(_2604_),
    .A2(_2607_),
    .ZN(_2636_));
 AOI21_X1 _3472_ (.A(_2636_),
    .B1(_2608_),
    .B2(_2565_),
    .ZN(_2637_));
 XNOR2_X1 _3473_ (.A(\section_2.xn2[9] ),
    .B(\section_2.xn2[8] ),
    .ZN(_2638_));
 INV_X1 _3474_ (.A(_0031_),
    .ZN(_2639_));
 AOI22_X1 _3475_ (.A1(_2639_),
    .A2(_2602_),
    .B1(_2603_),
    .B2(\section_2.xn2[9] ),
    .ZN(_2640_));
 NAND3_X1 _3476_ (.A1(_2500_),
    .A2(_2531_),
    .A3(_2601_),
    .ZN(_2641_));
 AND2_X1 _3477_ (.A1(_2568_),
    .A2(_2600_),
    .ZN(_2642_));
 AOI21_X1 _3478_ (.A(_2642_),
    .B1(_2601_),
    .B2(_2566_),
    .ZN(_2643_));
 NAND2_X1 _3479_ (.A1(_2641_),
    .A2(_2643_),
    .ZN(_2644_));
 NOR2_X1 _3480_ (.A1(_2570_),
    .A2(_2599_),
    .ZN(_2645_));
 NOR3_X1 _3481_ (.A1(_0008_),
    .A2(_2524_),
    .A3(_2597_),
    .ZN(_2646_));
 AOI21_X1 _3482_ (.A(_2646_),
    .B1(_2598_),
    .B2(_0003_),
    .ZN(_2647_));
 NOR2_X1 _3483_ (.A1(_0030_),
    .A2(_2596_),
    .ZN(_2648_));
 NOR2_X1 _3484_ (.A1(_2578_),
    .A2(_2594_),
    .ZN(_2649_));
 AOI21_X1 _3485_ (.A(_2649_),
    .B1(_2595_),
    .B2(_2577_),
    .ZN(_2650_));
 AND2_X1 _3486_ (.A1(_2508_),
    .A2(_2519_),
    .ZN(_2651_));
 OAI21_X1 _3487_ (.A(_2593_),
    .B1(_2651_),
    .B2(_2579_),
    .ZN(_2652_));
 NOR2_X1 _3488_ (.A1(_2583_),
    .A2(_2591_),
    .ZN(_2653_));
 AOI21_X1 _3489_ (.A(_2653_),
    .B1(_2592_),
    .B2(_2581_),
    .ZN(_2654_));
 NAND2_X1 _3490_ (.A1(\coll_reg[7] ),
    .A2(\coll_reg[5] ),
    .ZN(_2655_));
 OR2_X1 _3491_ (.A1(_2587_),
    .A2(_2589_),
    .ZN(_2656_));
 OAI21_X1 _3492_ (.A(_2656_),
    .B1(_2590_),
    .B2(_2584_),
    .ZN(_2657_));
 XOR2_X1 _3493_ (.A(\coll_reg[8] ),
    .B(\coll_reg[6] ),
    .Z(_2658_));
 AND2_X1 _3494_ (.A1(\coll_reg[8] ),
    .A2(\coll_reg[10] ),
    .ZN(_2659_));
 OR2_X1 _3495_ (.A1(\coll_reg[9] ),
    .A2(_2659_),
    .ZN(_2660_));
 OAI21_X1 _3496_ (.A(\coll_reg[9] ),
    .B1(\coll_reg[8] ),
    .B2(\coll_reg[10] ),
    .ZN(_2661_));
 NAND2_X1 _3497_ (.A1(_2660_),
    .A2(_2661_),
    .ZN(_2662_));
 XNOR2_X1 _3498_ (.A(_2658_),
    .B(_2662_),
    .ZN(_2663_));
 XNOR2_X1 _3499_ (.A(_2657_),
    .B(_2663_),
    .ZN(_2664_));
 XOR2_X1 _3500_ (.A(_2655_),
    .B(_2664_),
    .Z(_2665_));
 XOR2_X1 _3501_ (.A(_2654_),
    .B(_2665_),
    .Z(_2666_));
 XOR2_X1 _3502_ (.A(_2652_),
    .B(_2666_),
    .Z(_2667_));
 XNOR2_X1 _3503_ (.A(_2650_),
    .B(_2667_),
    .ZN(_2668_));
 XNOR2_X1 _3504_ (.A(\section_1.yn2[10] ),
    .B(_2668_),
    .ZN(_2669_));
 XNOR2_X1 _3505_ (.A(_2648_),
    .B(_2669_),
    .ZN(_2670_));
 XNOR2_X1 _3506_ (.A(_2443_),
    .B(_2670_),
    .ZN(_2671_));
 XNOR2_X1 _3507_ (.A(_2647_),
    .B(_2671_),
    .ZN(_2672_));
 XNOR2_X1 _3508_ (.A(_2645_),
    .B(_2672_),
    .ZN(_2673_));
 XNOR2_X1 _3509_ (.A(_2644_),
    .B(_2673_),
    .ZN(_2674_));
 XNOR2_X1 _3510_ (.A(_2640_),
    .B(_2674_),
    .ZN(_2675_));
 XNOR2_X1 _3511_ (.A(_2638_),
    .B(_2675_),
    .ZN(_2676_));
 XOR2_X1 _3512_ (.A(_2637_),
    .B(_2676_),
    .Z(_2677_));
 XNOR2_X1 _3513_ (.A(_2635_),
    .B(_2677_),
    .ZN(_2678_));
 XOR2_X1 _3514_ (.A(_2633_),
    .B(_2678_),
    .Z(_2679_));
 XNOR2_X1 _3515_ (.A(_2631_),
    .B(_2679_),
    .ZN(_2680_));
 XOR2_X1 _3516_ (.A(_2630_),
    .B(_2680_),
    .Z(_2681_));
 XNOR2_X1 _3517_ (.A(_2628_),
    .B(_2681_),
    .ZN(_2682_));
 XNOR2_X1 _3518_ (.A(_2626_),
    .B(_2682_),
    .ZN(_2683_));
 XOR2_X1 _3519_ (.A(_2625_),
    .B(_2683_),
    .Z(_2684_));
 XOR2_X1 _3520_ (.A(_2624_),
    .B(_2684_),
    .Z(_2685_));
 XNOR2_X1 _3521_ (.A(_2623_),
    .B(_2685_),
    .ZN(_2686_));
 NOR2_X1 _3522_ (.A1(_2620_),
    .A2(_2686_),
    .ZN(_2687_));
 NOR2_X1 _3523_ (.A1(z[2]),
    .A2(_2621_),
    .ZN(_2688_));
 NAND2_X1 _3524_ (.A1(_2624_),
    .A2(_2684_),
    .ZN(_2689_));
 NOR2_X1 _3525_ (.A1(_2624_),
    .A2(_2684_),
    .ZN(_2690_));
 INV_X1 _3526_ (.A(_2623_),
    .ZN(_2691_));
 OAI21_X1 _3527_ (.A(_2689_),
    .B1(_2690_),
    .B2(_2691_),
    .ZN(_2692_));
 NAND2_X1 _3528_ (.A1(z[2]),
    .A2(z[1]),
    .ZN(_2693_));
 XOR2_X1 _3529_ (.A(z[3]),
    .B(z[2]),
    .Z(_2694_));
 XNOR2_X1 _3530_ (.A(_2693_),
    .B(_2694_),
    .ZN(_2695_));
 INV_X1 _3531_ (.A(_2695_),
    .ZN(_2696_));
 NAND2_X1 _3532_ (.A1(_2625_),
    .A2(_2683_),
    .ZN(_2697_));
 NAND2_X1 _3533_ (.A1(z[8]),
    .A2(_2682_),
    .ZN(_2698_));
 NOR2_X1 _3534_ (.A1(_2630_),
    .A2(_2680_),
    .ZN(_2699_));
 AOI21_X1 _3535_ (.A(_2699_),
    .B1(_2681_),
    .B2(_2627_),
    .ZN(_2700_));
 NAND3_X1 _3536_ (.A1(_2554_),
    .A2(_2614_),
    .A3(_2681_),
    .ZN(_2701_));
 NOR2_X1 _3537_ (.A1(_2633_),
    .A2(_2678_),
    .ZN(_2702_));
 AOI21_X1 _3538_ (.A(_2702_),
    .B1(_2679_),
    .B2(_2631_),
    .ZN(_2703_));
 NOR2_X1 _3539_ (.A1(_0020_),
    .A2(_2634_),
    .ZN(_2704_));
 NOR2_X1 _3540_ (.A1(_2637_),
    .A2(_2676_),
    .ZN(_2705_));
 AOI21_X1 _3541_ (.A(_2705_),
    .B1(_2677_),
    .B2(_2635_),
    .ZN(_2706_));
 NAND2_X1 _3542_ (.A1(\section_2.xn2[9] ),
    .A2(\section_2.xn2[8] ),
    .ZN(_2707_));
 XOR2_X1 _3543_ (.A(_0018_),
    .B(_2707_),
    .Z(_2708_));
 OR2_X1 _3544_ (.A1(_2640_),
    .A2(_2674_),
    .ZN(_2709_));
 OAI21_X1 _3545_ (.A(_2709_),
    .B1(_2675_),
    .B2(_2638_),
    .ZN(_2710_));
 XOR2_X1 _3546_ (.A(\section_2.xn2[10] ),
    .B(\section_2.xn2[9] ),
    .Z(_2711_));
 INV_X1 _3547_ (.A(_2645_),
    .ZN(_2712_));
 NOR2_X1 _3548_ (.A1(_2712_),
    .A2(_2672_),
    .ZN(_2713_));
 AND2_X1 _3549_ (.A1(_2712_),
    .A2(_2672_),
    .ZN(_2714_));
 AOI211_X1 _3550_ (.A(_2713_),
    .B(_2714_),
    .C1(_2641_),
    .C2(_2643_),
    .ZN(_2715_));
 NOR2_X1 _3551_ (.A1(_2647_),
    .A2(_2671_),
    .ZN(_2716_));
 INV_X1 _3552_ (.A(\section_1.yn2[10] ),
    .ZN(_2717_));
 NOR2_X1 _3553_ (.A1(_2717_),
    .A2(_2668_),
    .ZN(_2718_));
 NOR2_X1 _3554_ (.A1(_2652_),
    .A2(_2666_),
    .ZN(_2719_));
 AOI21_X1 _3555_ (.A(_2719_),
    .B1(_2667_),
    .B2(_2649_),
    .ZN(_2720_));
 NAND2_X1 _3556_ (.A1(_2595_),
    .A2(_2667_),
    .ZN(_2721_));
 OR2_X1 _3557_ (.A1(_2576_),
    .A2(_2721_),
    .ZN(_2722_));
 OAI221_X1 _3558_ (.A(_2720_),
    .B1(_2721_),
    .B2(_2575_),
    .C1(_2464_),
    .C2(_2722_),
    .ZN(_2723_));
 INV_X1 _3559_ (.A(_2665_),
    .ZN(_2724_));
 NOR2_X1 _3560_ (.A1(_2654_),
    .A2(_2724_),
    .ZN(_2725_));
 NOR2_X1 _3561_ (.A1(_2655_),
    .A2(_2664_),
    .ZN(_2726_));
 AOI21_X1 _3562_ (.A(_2726_),
    .B1(_2663_),
    .B2(_2657_),
    .ZN(_2727_));
 NAND2_X1 _3563_ (.A1(\coll_reg[8] ),
    .A2(\coll_reg[6] ),
    .ZN(_2728_));
 XOR2_X1 _3564_ (.A(\coll_reg[9] ),
    .B(\coll_reg[7] ),
    .Z(_2729_));
 NAND3_X1 _3565_ (.A1(_2658_),
    .A2(_2660_),
    .A3(_2661_),
    .ZN(_2730_));
 NAND2_X1 _3566_ (.A1(\coll_reg[9] ),
    .A2(\coll_reg[10] ),
    .ZN(_2731_));
 NAND2_X1 _3567_ (.A1(\coll_reg[8] ),
    .A2(\coll_reg[10] ),
    .ZN(_2732_));
 NAND2_X1 _3568_ (.A1(_2731_),
    .A2(_2732_),
    .ZN(_2733_));
 NOR2_X1 _3569_ (.A1(_2588_),
    .A2(_2733_),
    .ZN(_2734_));
 OAI21_X1 _3570_ (.A(_2730_),
    .B1(_2734_),
    .B2(_0000_),
    .ZN(_2735_));
 XOR2_X1 _3571_ (.A(_2729_),
    .B(_2735_),
    .Z(_2736_));
 XNOR2_X1 _3572_ (.A(_2728_),
    .B(_2736_),
    .ZN(_2737_));
 XNOR2_X1 _3573_ (.A(_2727_),
    .B(_2737_),
    .ZN(_2738_));
 XNOR2_X1 _3574_ (.A(_2725_),
    .B(_2738_),
    .ZN(_2739_));
 XNOR2_X1 _3575_ (.A(_2723_),
    .B(_2739_),
    .ZN(_2740_));
 XOR2_X1 _3576_ (.A(_2718_),
    .B(_2740_),
    .Z(_2741_));
 XOR2_X1 _3577_ (.A(_0008_),
    .B(_2741_),
    .Z(_2742_));
 NOR3_X1 _3578_ (.A1(_0030_),
    .A2(_2596_),
    .A3(_2669_),
    .ZN(_2743_));
 AOI21_X1 _3579_ (.A(_2743_),
    .B1(_2670_),
    .B2(_0001_),
    .ZN(_2744_));
 XNOR2_X1 _3580_ (.A(_2742_),
    .B(_2744_),
    .ZN(_2745_));
 XOR2_X1 _3581_ (.A(_2716_),
    .B(_2745_),
    .Z(_2746_));
 OR3_X1 _3582_ (.A1(_2713_),
    .A2(_2715_),
    .A3(_2746_),
    .ZN(_2747_));
 OAI21_X1 _3583_ (.A(_2746_),
    .B1(_2715_),
    .B2(_2713_),
    .ZN(_2748_));
 AND3_X1 _3584_ (.A1(_2639_),
    .A2(_2747_),
    .A3(_2748_),
    .ZN(_2749_));
 AOI21_X1 _3585_ (.A(_2639_),
    .B1(_2747_),
    .B2(_2748_),
    .ZN(_2750_));
 NOR2_X1 _3586_ (.A1(_2749_),
    .A2(_2750_),
    .ZN(_2751_));
 XOR2_X1 _3587_ (.A(_2711_),
    .B(_2751_),
    .Z(_2752_));
 XOR2_X1 _3588_ (.A(_2710_),
    .B(_2752_),
    .Z(_2753_));
 XNOR2_X1 _3589_ (.A(_2708_),
    .B(_2753_),
    .ZN(_2754_));
 XOR2_X1 _3590_ (.A(_2706_),
    .B(_2754_),
    .Z(_2755_));
 XNOR2_X1 _3591_ (.A(_2704_),
    .B(_2755_),
    .ZN(_2756_));
 XOR2_X1 _3592_ (.A(_2703_),
    .B(_2756_),
    .Z(_2757_));
 INV_X1 _3593_ (.A(_2757_),
    .ZN(_2758_));
 NAND3_X1 _3594_ (.A1(_2700_),
    .A2(_2701_),
    .A3(_2758_),
    .ZN(_2759_));
 AND3_X1 _3595_ (.A1(_2554_),
    .A2(_2614_),
    .A3(_2681_),
    .ZN(_2760_));
 OR2_X1 _3596_ (.A1(_2630_),
    .A2(_2680_),
    .ZN(_2761_));
 AND2_X1 _3597_ (.A1(_2630_),
    .A2(_2680_),
    .ZN(_2762_));
 OR2_X1 _3598_ (.A1(_2557_),
    .A2(_2613_),
    .ZN(_2763_));
 OAI21_X1 _3599_ (.A(_2761_),
    .B1(_2762_),
    .B2(_2763_),
    .ZN(_2764_));
 OAI21_X1 _3600_ (.A(_2757_),
    .B1(_2760_),
    .B2(_2764_),
    .ZN(_2765_));
 AOI21_X1 _3601_ (.A(z[9]),
    .B1(_2759_),
    .B2(_2765_),
    .ZN(_2766_));
 INV_X1 _3602_ (.A(net69),
    .ZN(_2767_));
 NOR3_X1 _3603_ (.A1(_2764_),
    .A2(_2760_),
    .A3(_2757_),
    .ZN(_2768_));
 AOI21_X1 _3604_ (.A(_2758_),
    .B1(_2701_),
    .B2(_2700_),
    .ZN(_2769_));
 NOR3_X1 _3605_ (.A1(_2767_),
    .A2(_2768_),
    .A3(_2769_),
    .ZN(_2770_));
 NOR3_X1 _3606_ (.A1(_2698_),
    .A2(_2766_),
    .A3(_2770_),
    .ZN(_2771_));
 AND2_X1 _3607_ (.A1(z[8]),
    .A2(_2682_),
    .ZN(_2772_));
 OAI21_X1 _3608_ (.A(_2767_),
    .B1(_2768_),
    .B2(_2769_),
    .ZN(_2773_));
 NAND3_X1 _3609_ (.A1(z[9]),
    .A2(_2759_),
    .A3(_2765_),
    .ZN(_2774_));
 AOI21_X1 _3610_ (.A(_2772_),
    .B1(_2773_),
    .B2(_2774_),
    .ZN(_2775_));
 NOR3_X1 _3611_ (.A1(_2697_),
    .A2(_2771_),
    .A3(_2775_),
    .ZN(_2776_));
 NAND3_X1 _3612_ (.A1(_2772_),
    .A2(_2773_),
    .A3(_2774_),
    .ZN(_2777_));
 OAI21_X1 _3613_ (.A(_2698_),
    .B1(_2766_),
    .B2(_2770_),
    .ZN(_2778_));
 AOI22_X1 _3614_ (.A1(_2625_),
    .A2(_2683_),
    .B1(_2777_),
    .B2(_2778_),
    .ZN(_2779_));
 OAI21_X1 _3615_ (.A(_2696_),
    .B1(_2776_),
    .B2(_2779_),
    .ZN(_2780_));
 OR3_X1 _3616_ (.A1(_2697_),
    .A2(_2771_),
    .A3(_2775_),
    .ZN(_2781_));
 OAI21_X1 _3617_ (.A(_2697_),
    .B1(_2771_),
    .B2(_2775_),
    .ZN(_2782_));
 NAND3_X1 _3618_ (.A1(_2695_),
    .A2(_2781_),
    .A3(_2782_),
    .ZN(_2783_));
 NAND3_X1 _3619_ (.A1(_2692_),
    .A2(_2780_),
    .A3(_2783_),
    .ZN(_2784_));
 AOI22_X1 _3620_ (.A1(_2624_),
    .A2(_2684_),
    .B1(_2685_),
    .B2(_2623_),
    .ZN(_2785_));
 AOI21_X1 _3621_ (.A(_2695_),
    .B1(_2781_),
    .B2(_2782_),
    .ZN(_2786_));
 NOR3_X1 _3622_ (.A1(_2696_),
    .A2(_2776_),
    .A3(_2779_),
    .ZN(_2787_));
 OAI21_X1 _3623_ (.A(_2785_),
    .B1(_2786_),
    .B2(_2787_),
    .ZN(_2788_));
 NAND3_X1 _3624_ (.A1(_2688_),
    .A2(_2784_),
    .A3(_2788_),
    .ZN(_2789_));
 OR2_X1 _3625_ (.A1(z[2]),
    .A2(_2621_),
    .ZN(_2790_));
 NOR3_X1 _3626_ (.A1(_2785_),
    .A2(_2786_),
    .A3(_2787_),
    .ZN(_2791_));
 AOI21_X1 _3627_ (.A(_2692_),
    .B1(_2780_),
    .B2(_2783_),
    .ZN(_2792_));
 OAI21_X1 _3628_ (.A(_2790_),
    .B1(_2791_),
    .B2(_2792_),
    .ZN(_2793_));
 NAND3_X1 _3629_ (.A1(_2687_),
    .A2(_2789_),
    .A3(_2793_),
    .ZN(_2794_));
 NAND2_X1 _3630_ (.A1(_2784_),
    .A2(_2789_),
    .ZN(_2795_));
 OR2_X1 _3631_ (.A1(z[3]),
    .A2(_2693_),
    .ZN(_2796_));
 NAND2_X1 _3632_ (.A1(_2781_),
    .A2(_2783_),
    .ZN(_2797_));
 NAND2_X1 _3633_ (.A1(z[3]),
    .A2(z[2]),
    .ZN(_2798_));
 XOR2_X1 _3634_ (.A(z[4]),
    .B(z[3]),
    .Z(_2799_));
 XNOR2_X1 _3635_ (.A(_2798_),
    .B(_2799_),
    .ZN(_2800_));
 NOR2_X1 _3636_ (.A1(_2706_),
    .A2(_2754_),
    .ZN(_2801_));
 AOI21_X1 _3637_ (.A(_2801_),
    .B1(_2755_),
    .B2(_2704_),
    .ZN(_2802_));
 OR2_X1 _3638_ (.A1(_0018_),
    .A2(_2707_),
    .ZN(_2803_));
 AND2_X1 _3639_ (.A1(_2710_),
    .A2(_2752_),
    .ZN(_2804_));
 AOI21_X1 _3640_ (.A(_2804_),
    .B1(_2753_),
    .B2(_2708_),
    .ZN(_2805_));
 NAND2_X1 _3641_ (.A1(\section_2.xn2[10] ),
    .A2(\section_2.xn2[9] ),
    .ZN(_2806_));
 XOR2_X1 _3642_ (.A(_0016_),
    .B(_2806_),
    .Z(_2807_));
 AOI21_X1 _3643_ (.A(_2749_),
    .B1(_2751_),
    .B2(_2711_),
    .ZN(_2808_));
 NOR2_X1 _3644_ (.A1(_2568_),
    .A2(_2600_),
    .ZN(_2809_));
 NAND2_X1 _3645_ (.A1(_2568_),
    .A2(_2600_),
    .ZN(_2810_));
 OR2_X1 _3646_ (.A1(_2502_),
    .A2(_2530_),
    .ZN(_2811_));
 AOI21_X1 _3647_ (.A(_2809_),
    .B1(_2810_),
    .B2(_2811_),
    .ZN(_2812_));
 NAND3_X1 _3648_ (.A1(_2812_),
    .A2(_2673_),
    .A3(_2746_),
    .ZN(_2813_));
 AND2_X1 _3649_ (.A1(_2716_),
    .A2(_2745_),
    .ZN(_2814_));
 AOI21_X1 _3650_ (.A(_2814_),
    .B1(_2746_),
    .B2(_2713_),
    .ZN(_2815_));
 INV_X1 _3651_ (.A(_2500_),
    .ZN(_2816_));
 NAND4_X1 _3652_ (.A1(_2531_),
    .A2(_2601_),
    .A3(_2673_),
    .A4(_2746_),
    .ZN(_2817_));
 OAI211_X1 _3653_ (.A(_2813_),
    .B(_2815_),
    .C1(_2816_),
    .C2(_2817_),
    .ZN(_2818_));
 INV_X1 _3654_ (.A(_2742_),
    .ZN(_2819_));
 NOR2_X1 _3655_ (.A1(_2819_),
    .A2(_2744_),
    .ZN(_2820_));
 NOR2_X1 _3656_ (.A1(_2717_),
    .A2(_2740_),
    .ZN(_2821_));
 AOI22_X1 _3657_ (.A1(_2668_),
    .A2(_2821_),
    .B1(_2741_),
    .B2(_0008_),
    .ZN(_2822_));
 INV_X1 _3658_ (.A(_2737_),
    .ZN(_2823_));
 NOR2_X1 _3659_ (.A1(_2727_),
    .A2(_2823_),
    .ZN(_2824_));
 NAND2_X1 _3660_ (.A1(_2729_),
    .A2(_2735_),
    .ZN(_2825_));
 NOR2_X1 _3661_ (.A1(_2729_),
    .A2(_2735_),
    .ZN(_2826_));
 OAI21_X1 _3662_ (.A(_2825_),
    .B1(_2826_),
    .B2(_2728_),
    .ZN(_2827_));
 AOI21_X1 _3663_ (.A(\coll_reg[8] ),
    .B1(\coll_reg[7] ),
    .B2(\coll_reg[9] ),
    .ZN(_2828_));
 AOI21_X1 _3664_ (.A(_2828_),
    .B1(_2588_),
    .B2(\coll_reg[7] ),
    .ZN(_2829_));
 XOR2_X1 _3665_ (.A(_2827_),
    .B(_2829_),
    .Z(_2830_));
 XOR2_X1 _3666_ (.A(_2824_),
    .B(_2830_),
    .Z(_2831_));
 AND2_X1 _3667_ (.A1(_2725_),
    .A2(_2738_),
    .ZN(_2832_));
 INV_X1 _3668_ (.A(_2739_),
    .ZN(_2833_));
 AOI21_X1 _3669_ (.A(_2832_),
    .B1(_2833_),
    .B2(_2723_),
    .ZN(_2834_));
 XNOR2_X1 _3670_ (.A(_2831_),
    .B(_2834_),
    .ZN(_2835_));
 XOR2_X1 _3671_ (.A(_2821_),
    .B(_2835_),
    .Z(_2836_));
 XOR2_X1 _3672_ (.A(_0030_),
    .B(_2836_),
    .Z(_2837_));
 XNOR2_X1 _3673_ (.A(_2822_),
    .B(_2837_),
    .ZN(_2838_));
 XNOR2_X1 _3674_ (.A(_2820_),
    .B(_2838_),
    .ZN(_2839_));
 XNOR2_X1 _3675_ (.A(_2818_),
    .B(_2839_),
    .ZN(_2840_));
 XNOR2_X1 _3676_ (.A(\section_2.xn2[10] ),
    .B(_2840_),
    .ZN(_2841_));
 XNOR2_X1 _3677_ (.A(_2808_),
    .B(_2841_),
    .ZN(_2842_));
 XOR2_X1 _3678_ (.A(_2807_),
    .B(_2842_),
    .Z(_2843_));
 XNOR2_X1 _3679_ (.A(_2805_),
    .B(_2843_),
    .ZN(_2844_));
 XNOR2_X1 _3680_ (.A(_2803_),
    .B(_2844_),
    .ZN(_2845_));
 XOR2_X1 _3681_ (.A(_2802_),
    .B(_2845_),
    .Z(_2846_));
 NAND2_X1 _3682_ (.A1(_2757_),
    .A2(_2846_),
    .ZN(_2847_));
 AOI21_X1 _3683_ (.A(_2847_),
    .B1(_2701_),
    .B2(_2700_),
    .ZN(_2848_));
 NOR2_X1 _3684_ (.A1(_2703_),
    .A2(_2756_),
    .ZN(_2849_));
 NAND2_X1 _3685_ (.A1(_2849_),
    .A2(_2846_),
    .ZN(_2850_));
 INV_X1 _3686_ (.A(_2850_),
    .ZN(_2851_));
 NOR2_X1 _3687_ (.A1(_2849_),
    .A2(_2846_),
    .ZN(_2852_));
 AOI211_X1 _3688_ (.A(_2848_),
    .B(_2851_),
    .C1(_2765_),
    .C2(_2852_),
    .ZN(_2853_));
 XNOR2_X1 _3689_ (.A(z[10]),
    .B(_2853_),
    .ZN(_2854_));
 XNOR2_X1 _3690_ (.A(_2774_),
    .B(_2854_),
    .ZN(_2855_));
 XNOR2_X1 _3691_ (.A(_2777_),
    .B(_2855_),
    .ZN(_2856_));
 XNOR2_X1 _3692_ (.A(_2800_),
    .B(_2856_),
    .ZN(_2857_));
 XNOR2_X1 _3693_ (.A(_2797_),
    .B(_2857_),
    .ZN(_2858_));
 XOR2_X1 _3694_ (.A(_2796_),
    .B(_2858_),
    .Z(_2859_));
 XNOR2_X1 _3695_ (.A(_2795_),
    .B(_2859_),
    .ZN(_2860_));
 XNOR2_X1 _3696_ (.A(_2794_),
    .B(_2860_),
    .ZN(_2861_));
 INV_X1 _3697_ (.A(net60),
    .ZN(_2862_));
 XOR2_X1 _3698_ (.A(_2374_),
    .B(_2424_),
    .Z(_2863_));
 NAND2_X1 _3699_ (.A1(z[4]),
    .A2(_2863_),
    .ZN(_2864_));
 XNOR2_X1 _3700_ (.A(z[5]),
    .B(_2486_),
    .ZN(_2865_));
 NOR2_X1 _3701_ (.A1(_2864_),
    .A2(_2865_),
    .ZN(_2866_));
 XOR2_X1 _3702_ (.A(_2487_),
    .B(_2548_),
    .Z(_2867_));
 XNOR2_X1 _3703_ (.A(_2866_),
    .B(_2867_),
    .ZN(_2868_));
 NOR2_X1 _3704_ (.A1(_2862_),
    .A2(_2868_),
    .ZN(_2869_));
 AOI21_X1 _3705_ (.A(_2869_),
    .B1(_2867_),
    .B2(_2866_),
    .ZN(_2870_));
 XNOR2_X1 _3706_ (.A(_1275_),
    .B(_2618_),
    .ZN(_2871_));
 NOR2_X1 _3707_ (.A1(_2870_),
    .A2(_2871_),
    .ZN(_2872_));
 XOR2_X1 _3708_ (.A(_2620_),
    .B(_2686_),
    .Z(_2873_));
 NAND2_X1 _3709_ (.A1(_2872_),
    .A2(_2873_),
    .ZN(_2874_));
 AOI21_X1 _3710_ (.A(_2687_),
    .B1(_2789_),
    .B2(_2793_),
    .ZN(_2875_));
 INV_X1 _3711_ (.A(_2687_),
    .ZN(_2876_));
 NOR3_X1 _3712_ (.A1(_2790_),
    .A2(_2791_),
    .A3(_2792_),
    .ZN(_2877_));
 AOI21_X1 _3713_ (.A(_2688_),
    .B1(_2784_),
    .B2(_2788_),
    .ZN(_2878_));
 NOR3_X1 _3714_ (.A1(_2876_),
    .A2(_2877_),
    .A3(_2878_),
    .ZN(_2879_));
 OAI21_X1 _3715_ (.A(_2874_),
    .B1(_2875_),
    .B2(_2879_),
    .ZN(_2880_));
 NOR3_X1 _3716_ (.A1(_2879_),
    .A2(_2874_),
    .A3(_2875_),
    .ZN(_2881_));
 XOR2_X1 _3717_ (.A(_2418_),
    .B(_2421_),
    .Z(_2882_));
 NAND2_X1 _3718_ (.A1(z[3]),
    .A2(_2882_),
    .ZN(_2883_));
 XNOR2_X1 _3719_ (.A(z[4]),
    .B(_2863_),
    .ZN(_2884_));
 NOR2_X1 _3720_ (.A1(_2883_),
    .A2(_2884_),
    .ZN(_2885_));
 XOR2_X1 _3721_ (.A(_2864_),
    .B(_2865_),
    .Z(_2886_));
 AND2_X1 _3722_ (.A1(_2885_),
    .A2(_2886_),
    .ZN(_2887_));
 INV_X1 _3723_ (.A(_2887_),
    .ZN(_2888_));
 XNOR2_X1 _3724_ (.A(_2862_),
    .B(_2868_),
    .ZN(_2889_));
 NOR2_X1 _3725_ (.A1(_2888_),
    .A2(_2889_),
    .ZN(_2890_));
 XOR2_X1 _3726_ (.A(_2870_),
    .B(_2871_),
    .Z(_2891_));
 NAND2_X1 _3727_ (.A1(_2890_),
    .A2(_2891_),
    .ZN(_2892_));
 XNOR2_X1 _3728_ (.A(_2872_),
    .B(_2873_),
    .ZN(_2893_));
 OR2_X1 _3729_ (.A1(_2892_),
    .A2(_2893_),
    .ZN(_2894_));
 XNOR2_X1 _3730_ (.A(_2414_),
    .B(_2416_),
    .ZN(_2895_));
 NAND2_X1 _3731_ (.A1(z[2]),
    .A2(_2895_),
    .ZN(_2896_));
 XNOR2_X1 _3732_ (.A(z[3]),
    .B(_2882_),
    .ZN(_2897_));
 NOR2_X1 _3733_ (.A1(_2896_),
    .A2(_2897_),
    .ZN(_2898_));
 XOR2_X1 _3734_ (.A(_2883_),
    .B(_2884_),
    .Z(_2899_));
 AND2_X1 _3735_ (.A1(_2898_),
    .A2(_2899_),
    .ZN(_2900_));
 XNOR2_X1 _3736_ (.A(_2887_),
    .B(_2889_),
    .ZN(_2901_));
 AND3_X1 _3737_ (.A1(_2886_),
    .A2(_2900_),
    .A3(_2901_),
    .ZN(_2902_));
 NOR2_X1 _3738_ (.A1(_2890_),
    .A2(_2902_),
    .ZN(_2903_));
 XNOR2_X1 _3739_ (.A(_2891_),
    .B(_2903_),
    .ZN(_2904_));
 NAND2_X1 _3740_ (.A1(_2886_),
    .A2(_2900_),
    .ZN(_2905_));
 XNOR2_X1 _3741_ (.A(_2905_),
    .B(_2901_),
    .ZN(_2906_));
 XOR2_X1 _3742_ (.A(_2412_),
    .B(_2413_),
    .Z(_2907_));
 NAND2_X1 _3743_ (.A1(z[1]),
    .A2(_2907_),
    .ZN(_2908_));
 XNOR2_X1 _3744_ (.A(z[2]),
    .B(_2895_),
    .ZN(_2909_));
 NOR2_X1 _3745_ (.A1(_2908_),
    .A2(_2909_),
    .ZN(_2910_));
 XOR2_X1 _3746_ (.A(_2896_),
    .B(_2897_),
    .Z(_2911_));
 AND2_X1 _3747_ (.A1(_2910_),
    .A2(_2911_),
    .ZN(_2912_));
 XOR2_X1 _3748_ (.A(_2898_),
    .B(_2899_),
    .Z(_2913_));
 NAND2_X1 _3749_ (.A1(_2912_),
    .A2(_2913_),
    .ZN(_2914_));
 NOR2_X1 _3750_ (.A1(_2885_),
    .A2(_2900_),
    .ZN(_2915_));
 XOR2_X1 _3751_ (.A(_2886_),
    .B(_2915_),
    .Z(_2916_));
 NOR2_X1 _3752_ (.A1(_2914_),
    .A2(_2916_),
    .ZN(_2917_));
 NAND2_X1 _3753_ (.A1(_2906_),
    .A2(_2917_),
    .ZN(_2918_));
 XNOR2_X1 _3754_ (.A(_2410_),
    .B(_2411_),
    .ZN(_2919_));
 OR2_X1 _3755_ (.A1(_2862_),
    .A2(_2919_),
    .ZN(_2920_));
 XNOR2_X1 _3756_ (.A(z[1]),
    .B(_2907_),
    .ZN(_2921_));
 NOR2_X1 _3757_ (.A1(_2920_),
    .A2(_2921_),
    .ZN(_2922_));
 XOR2_X1 _3758_ (.A(_2908_),
    .B(_2909_),
    .Z(_2923_));
 AND2_X1 _3759_ (.A1(_2922_),
    .A2(_2923_),
    .ZN(_2924_));
 XOR2_X1 _3760_ (.A(_2910_),
    .B(_2911_),
    .Z(_2925_));
 NAND2_X1 _3761_ (.A1(_2924_),
    .A2(_2925_),
    .ZN(_2926_));
 XNOR2_X1 _3762_ (.A(_2912_),
    .B(_2913_),
    .ZN(_2927_));
 OR3_X1 _3763_ (.A1(_2916_),
    .A2(_2926_),
    .A3(_2927_),
    .ZN(_2928_));
 XNOR2_X1 _3764_ (.A(_2906_),
    .B(_2917_),
    .ZN(_2929_));
 OAI21_X1 _3765_ (.A(_2918_),
    .B1(_2928_),
    .B2(_2929_),
    .ZN(_2930_));
 AOI22_X1 _3766_ (.A1(_2891_),
    .A2(_2902_),
    .B1(_2904_),
    .B2(_2930_),
    .ZN(_2931_));
 XNOR2_X1 _3767_ (.A(_2892_),
    .B(_2893_),
    .ZN(_2932_));
 OAI21_X1 _3768_ (.A(_2894_),
    .B1(_2931_),
    .B2(_2932_),
    .ZN(_2933_));
 OAI21_X1 _3769_ (.A(_2880_),
    .B1(_2881_),
    .B2(_2933_),
    .ZN(_2934_));
 OAI22_X1 _3770_ (.A1(_2794_),
    .A2(_2860_),
    .B1(_2861_),
    .B2(_2934_),
    .ZN(_2935_));
 AND2_X1 _3771_ (.A1(_2795_),
    .A2(_2859_),
    .ZN(_2936_));
 NAND2_X1 _3772_ (.A1(_2797_),
    .A2(_2857_),
    .ZN(_2937_));
 OAI21_X1 _3773_ (.A(_2937_),
    .B1(_2858_),
    .B2(_2796_),
    .ZN(_2938_));
 NOR2_X1 _3774_ (.A1(z[4]),
    .A2(_2798_),
    .ZN(_2939_));
 INV_X1 _3775_ (.A(_2939_),
    .ZN(_2940_));
 NOR2_X1 _3776_ (.A1(_2777_),
    .A2(_2855_),
    .ZN(_2941_));
 NAND2_X1 _3777_ (.A1(_2777_),
    .A2(_2855_),
    .ZN(_2942_));
 AOI21_X1 _3778_ (.A(_2941_),
    .B1(_2942_),
    .B2(_2800_),
    .ZN(_2943_));
 NAND2_X1 _3779_ (.A1(z[4]),
    .A2(z[3]),
    .ZN(_2944_));
 NOR2_X1 _3780_ (.A1(z[5]),
    .A2(_2944_),
    .ZN(_2945_));
 OR2_X1 _3781_ (.A1(z[5]),
    .A2(z[4]),
    .ZN(_2946_));
 NAND2_X1 _3782_ (.A1(z[5]),
    .A2(z[4]),
    .ZN(_2947_));
 AOI22_X1 _3783_ (.A1(z[4]),
    .A2(z[3]),
    .B1(_2946_),
    .B2(_2947_),
    .ZN(_2948_));
 NOR2_X1 _3784_ (.A1(_2945_),
    .A2(_2948_),
    .ZN(_2949_));
 OR2_X1 _3785_ (.A1(_2774_),
    .A2(_2854_),
    .ZN(_2950_));
 INV_X1 _3786_ (.A(net81),
    .ZN(_2951_));
 NOR2_X1 _3787_ (.A1(_2951_),
    .A2(_2853_),
    .ZN(_2952_));
 OR2_X1 _3788_ (.A1(_2802_),
    .A2(_2845_),
    .ZN(_2953_));
 NAND2_X1 _3789_ (.A1(_2953_),
    .A2(_2850_),
    .ZN(_2954_));
 OR2_X1 _3790_ (.A1(_2805_),
    .A2(_2843_),
    .ZN(_2955_));
 AND2_X1 _3791_ (.A1(_2805_),
    .A2(_2843_),
    .ZN(_2956_));
 OAI21_X1 _3792_ (.A(_2955_),
    .B1(_2956_),
    .B2(_2803_),
    .ZN(_2957_));
 NOR2_X1 _3793_ (.A1(_0016_),
    .A2(_2806_),
    .ZN(_2958_));
 NOR2_X1 _3794_ (.A1(_2808_),
    .A2(_2841_),
    .ZN(_0120_));
 NAND2_X1 _3795_ (.A1(_2808_),
    .A2(_2841_),
    .ZN(_0121_));
 AOI21_X1 _3796_ (.A(_0120_),
    .B1(_0121_),
    .B2(_2807_),
    .ZN(_0122_));
 XOR2_X1 _3797_ (.A(\section_2.xn2[10] ),
    .B(_0031_),
    .Z(_0123_));
 XOR2_X1 _3798_ (.A(_2840_),
    .B(_0123_),
    .Z(_0124_));
 NOR2_X1 _3799_ (.A1(_0031_),
    .A2(_0124_),
    .ZN(_0125_));
 AND2_X1 _3800_ (.A1(_2820_),
    .A2(_2838_),
    .ZN(_0126_));
 INV_X1 _3801_ (.A(_2839_),
    .ZN(_0127_));
 AOI21_X1 _3802_ (.A(_0126_),
    .B1(_0127_),
    .B2(_2818_),
    .ZN(_0128_));
 INV_X1 _3803_ (.A(_2822_),
    .ZN(_0129_));
 NAND2_X1 _3804_ (.A1(_0129_),
    .A2(_2837_),
    .ZN(_0130_));
 NOR2_X1 _3805_ (.A1(_2717_),
    .A2(_2835_),
    .ZN(_0131_));
 NAND2_X1 _3806_ (.A1(_2740_),
    .A2(_0131_),
    .ZN(_0132_));
 NAND2_X1 _3807_ (.A1(_0030_),
    .A2(_2836_),
    .ZN(_0133_));
 AND2_X1 _3808_ (.A1(_2827_),
    .A2(_2829_),
    .ZN(_0134_));
 OAI21_X1 _3809_ (.A(_2660_),
    .B1(_2731_),
    .B2(_2585_),
    .ZN(_0135_));
 NAND2_X1 _3810_ (.A1(\coll_reg[7] ),
    .A2(_2588_),
    .ZN(_0136_));
 OAI21_X1 _3811_ (.A(_0136_),
    .B1(_0006_),
    .B2(\coll_reg[8] ),
    .ZN(_0137_));
 XNOR2_X1 _3812_ (.A(_0135_),
    .B(_0137_),
    .ZN(_0138_));
 XNOR2_X1 _3813_ (.A(_0134_),
    .B(_0138_),
    .ZN(_0139_));
 NOR2_X1 _3814_ (.A1(_2824_),
    .A2(_2830_),
    .ZN(_0140_));
 NAND2_X1 _3815_ (.A1(_2824_),
    .A2(_2830_),
    .ZN(_0141_));
 AOI21_X1 _3816_ (.A(_0140_),
    .B1(_2834_),
    .B2(_0141_),
    .ZN(_0142_));
 XNOR2_X1 _3817_ (.A(_0139_),
    .B(_0142_),
    .ZN(_0143_));
 INV_X1 _3818_ (.A(_0004_),
    .ZN(_0144_));
 XNOR2_X1 _3819_ (.A(_0144_),
    .B(_0131_),
    .ZN(_0145_));
 XNOR2_X1 _3820_ (.A(_0143_),
    .B(_0145_),
    .ZN(_0146_));
 AND3_X1 _3821_ (.A1(_0132_),
    .A2(_0133_),
    .A3(_0146_),
    .ZN(_0147_));
 AOI21_X1 _3822_ (.A(_0146_),
    .B1(_0133_),
    .B2(_0132_),
    .ZN(_0148_));
 OR2_X1 _3823_ (.A1(_0147_),
    .A2(_0148_),
    .ZN(_0149_));
 XNOR2_X1 _3824_ (.A(_0130_),
    .B(_0149_),
    .ZN(_0150_));
 XNOR2_X1 _3825_ (.A(_0123_),
    .B(_0150_),
    .ZN(_0151_));
 XNOR2_X1 _3826_ (.A(_0128_),
    .B(_0151_),
    .ZN(_0152_));
 XNOR2_X1 _3827_ (.A(_0031_),
    .B(_0152_),
    .ZN(_0153_));
 XNOR2_X1 _3828_ (.A(_0125_),
    .B(_0153_),
    .ZN(_0154_));
 XNOR2_X1 _3829_ (.A(_2711_),
    .B(_0154_),
    .ZN(_0155_));
 XOR2_X1 _3830_ (.A(_0122_),
    .B(_0155_),
    .Z(_0156_));
 XOR2_X1 _3831_ (.A(_2958_),
    .B(_0156_),
    .Z(_0157_));
 XOR2_X1 _3832_ (.A(_2957_),
    .B(_0157_),
    .Z(_0158_));
 OR3_X1 _3833_ (.A1(_2848_),
    .A2(_2954_),
    .A3(_0158_),
    .ZN(_0159_));
 OAI21_X1 _3834_ (.A(_0158_),
    .B1(_2954_),
    .B2(_2848_),
    .ZN(_0160_));
 AND2_X1 _3835_ (.A1(_0159_),
    .A2(_0160_),
    .ZN(_0161_));
 XNOR2_X1 _3836_ (.A(_2952_),
    .B(_0161_),
    .ZN(_0162_));
 XOR2_X1 _3837_ (.A(_2950_),
    .B(_0162_),
    .Z(_0163_));
 XNOR2_X1 _3838_ (.A(_2949_),
    .B(_0163_),
    .ZN(_0164_));
 XOR2_X1 _3839_ (.A(_2943_),
    .B(_0164_),
    .Z(_0165_));
 XNOR2_X1 _3840_ (.A(_2940_),
    .B(_0165_),
    .ZN(_0166_));
 XOR2_X1 _3841_ (.A(_2938_),
    .B(_0166_),
    .Z(_0167_));
 XNOR2_X1 _3842_ (.A(_2936_),
    .B(_0167_),
    .ZN(_0168_));
 XNOR2_X1 _3843_ (.A(_0002_),
    .B(\section_2.yn2[10] ),
    .ZN(_0169_));
 XNOR2_X1 _3844_ (.A(_0168_),
    .B(_0169_),
    .ZN(_0170_));
 XNOR2_X1 _3845_ (.A(_2935_),
    .B(_0170_),
    .ZN(_0171_));
 INV_X1 _3846_ (.A(_0171_),
    .ZN(_0172_));
 NOR2_X1 _3847_ (.A1(_0002_),
    .A2(_0172_),
    .ZN(_0173_));
 NAND2_X1 _3848_ (.A1(_2938_),
    .A2(_0166_),
    .ZN(_0174_));
 OR2_X1 _3849_ (.A1(_2943_),
    .A2(_0164_),
    .ZN(_0175_));
 AND2_X1 _3850_ (.A1(_2943_),
    .A2(_0164_),
    .ZN(_0176_));
 OAI21_X1 _3851_ (.A(_0175_),
    .B1(_0176_),
    .B2(_2940_),
    .ZN(_0177_));
 NOR2_X1 _3852_ (.A1(_2950_),
    .A2(_0162_),
    .ZN(_0178_));
 AOI21_X1 _3853_ (.A(_0178_),
    .B1(_0163_),
    .B2(_2949_),
    .ZN(_0179_));
 XOR2_X1 _3854_ (.A(z[6]),
    .B(z[5]),
    .Z(_0180_));
 XNOR2_X1 _3855_ (.A(_2947_),
    .B(_0180_),
    .ZN(_0181_));
 INV_X1 _3856_ (.A(_0181_),
    .ZN(_0182_));
 OR3_X1 _3857_ (.A1(_2951_),
    .A2(_2853_),
    .A3(_0161_),
    .ZN(_0183_));
 NAND2_X1 _3858_ (.A1(_2957_),
    .A2(_0157_),
    .ZN(_0184_));
 NOR2_X1 _3859_ (.A1(_0122_),
    .A2(_0155_),
    .ZN(_0185_));
 AOI21_X1 _3860_ (.A(_0185_),
    .B1(_0156_),
    .B2(_2958_),
    .ZN(_0186_));
 NAND2_X1 _3861_ (.A1(_2639_),
    .A2(_0152_),
    .ZN(_0187_));
 NOR2_X1 _3862_ (.A1(_0124_),
    .A2(_0187_),
    .ZN(_0188_));
 AOI21_X1 _3863_ (.A(_0188_),
    .B1(_0154_),
    .B2(_2711_),
    .ZN(_0189_));
 AND2_X1 _3864_ (.A1(_2717_),
    .A2(_0143_),
    .ZN(_0190_));
 NOR2_X1 _3865_ (.A1(_2717_),
    .A2(_0143_),
    .ZN(_0191_));
 AOI21_X1 _3866_ (.A(_0190_),
    .B1(_0191_),
    .B2(_2835_),
    .ZN(_0192_));
 INV_X1 _3867_ (.A(_0142_),
    .ZN(_0193_));
 NOR2_X1 _3868_ (.A1(_0139_),
    .A2(_0193_),
    .ZN(_0194_));
 AOI21_X1 _3869_ (.A(_0194_),
    .B1(_0138_),
    .B2(_0134_),
    .ZN(_0195_));
 NOR2_X1 _3870_ (.A1(_2585_),
    .A2(_2731_),
    .ZN(_0196_));
 AOI21_X1 _3871_ (.A(_0196_),
    .B1(_0137_),
    .B2(_2660_),
    .ZN(_0197_));
 NAND2_X1 _3872_ (.A1(_0195_),
    .A2(_0197_),
    .ZN(_0198_));
 XNOR2_X1 _3873_ (.A(_0004_),
    .B(_0191_),
    .ZN(_0199_));
 XNOR2_X1 _3874_ (.A(_0198_),
    .B(_0199_),
    .ZN(_0200_));
 XNOR2_X1 _3875_ (.A(_0192_),
    .B(_0200_),
    .ZN(_0201_));
 XNOR2_X1 _3876_ (.A(_0148_),
    .B(_0201_),
    .ZN(_0202_));
 OR2_X1 _3877_ (.A1(_0130_),
    .A2(_0149_),
    .ZN(_0203_));
 OAI21_X1 _3878_ (.A(_0203_),
    .B1(_0150_),
    .B2(_0128_),
    .ZN(_0204_));
 XOR2_X1 _3879_ (.A(_0202_),
    .B(_0204_),
    .Z(_0205_));
 XNOR2_X1 _3880_ (.A(_0187_),
    .B(_0205_),
    .ZN(_0206_));
 XOR2_X1 _3881_ (.A(_0189_),
    .B(_0206_),
    .Z(_0207_));
 XNOR2_X1 _3882_ (.A(_2806_),
    .B(_0207_),
    .ZN(_0208_));
 XNOR2_X1 _3883_ (.A(_0186_),
    .B(_0208_),
    .ZN(_0209_));
 INV_X1 _3884_ (.A(_0209_),
    .ZN(_0210_));
 AND3_X1 _3885_ (.A1(_0184_),
    .A2(_0160_),
    .A3(_0210_),
    .ZN(_0211_));
 AOI21_X1 _3886_ (.A(_0210_),
    .B1(_0160_),
    .B2(_0184_),
    .ZN(_0212_));
 OR2_X1 _3887_ (.A1(_0211_),
    .A2(_0212_),
    .ZN(_0213_));
 XNOR2_X1 _3888_ (.A(_0183_),
    .B(_0213_),
    .ZN(_0214_));
 XNOR2_X1 _3889_ (.A(_0182_),
    .B(_0214_),
    .ZN(_0215_));
 XOR2_X1 _3890_ (.A(_0179_),
    .B(_0215_),
    .Z(_0216_));
 XOR2_X1 _3891_ (.A(_2945_),
    .B(_0216_),
    .Z(_0217_));
 XNOR2_X1 _3892_ (.A(_0177_),
    .B(_0217_),
    .ZN(_0218_));
 XOR2_X1 _3893_ (.A(_0174_),
    .B(_0218_),
    .Z(_0219_));
 AND2_X1 _3894_ (.A1(_2936_),
    .A2(_0167_),
    .ZN(_0220_));
 OR2_X1 _3895_ (.A1(_2936_),
    .A2(_0167_),
    .ZN(_0221_));
 NOR2_X1 _3896_ (.A1(_2794_),
    .A2(_2860_),
    .ZN(_0222_));
 AOI21_X1 _3897_ (.A(_0220_),
    .B1(_0221_),
    .B2(_0222_),
    .ZN(_0223_));
 OR3_X1 _3898_ (.A1(_2861_),
    .A2(_2934_),
    .A3(_0168_),
    .ZN(_0224_));
 NAND2_X1 _3899_ (.A1(_0223_),
    .A2(_0224_),
    .ZN(_0225_));
 XNOR2_X1 _3900_ (.A(_0219_),
    .B(_0225_),
    .ZN(_0226_));
 XNOR2_X1 _3901_ (.A(_0169_),
    .B(_0226_),
    .ZN(_0227_));
 XOR2_X1 _3902_ (.A(_0173_),
    .B(_0227_),
    .Z(_0228_));
 NOR2_X1 _3903_ (.A1(_0002_),
    .A2(_0227_),
    .ZN(_0229_));
 AOI22_X1 _3904_ (.A1(_1264_),
    .A2(_0228_),
    .B1(_0229_),
    .B2(_0172_),
    .ZN(_0230_));
 XOR2_X1 _3905_ (.A(\section_2.yn2[10] ),
    .B(\section_2.yn2[9] ),
    .Z(_0231_));
 NOR2_X1 _3906_ (.A1(_0174_),
    .A2(_0218_),
    .ZN(_0232_));
 AOI21_X1 _3907_ (.A(_0232_),
    .B1(_0219_),
    .B2(_0225_),
    .ZN(_0233_));
 NAND2_X1 _3908_ (.A1(_0177_),
    .A2(_0217_),
    .ZN(_0234_));
 NOR2_X1 _3909_ (.A1(_0179_),
    .A2(_0215_),
    .ZN(_0235_));
 AOI21_X1 _3910_ (.A(_0235_),
    .B1(_0216_),
    .B2(_2945_),
    .ZN(_0236_));
 NOR2_X1 _3911_ (.A1(z[6]),
    .A2(_2947_),
    .ZN(_0237_));
 NAND3_X1 _3912_ (.A1(z[10]),
    .A2(_2853_),
    .A3(_0213_),
    .ZN(_0238_));
 OAI22_X1 _3913_ (.A1(_0182_),
    .A2(_0214_),
    .B1(_0238_),
    .B2(_0161_),
    .ZN(_0239_));
 NAND2_X1 _3914_ (.A1(z[6]),
    .A2(z[5]),
    .ZN(_0240_));
 NOR2_X1 _3915_ (.A1(z[7]),
    .A2(_0240_),
    .ZN(_0241_));
 OR2_X1 _3916_ (.A1(z[7]),
    .A2(z[6]),
    .ZN(_0242_));
 NAND2_X1 _3917_ (.A1(z[7]),
    .A2(z[6]),
    .ZN(_0243_));
 AOI22_X1 _3918_ (.A1(z[6]),
    .A2(z[5]),
    .B1(_0242_),
    .B2(_0243_),
    .ZN(_0244_));
 NOR2_X1 _3919_ (.A1(_0241_),
    .A2(_0244_),
    .ZN(_0245_));
 AOI21_X1 _3920_ (.A(_2951_),
    .B1(_0159_),
    .B2(_0160_),
    .ZN(_0246_));
 OAI21_X1 _3921_ (.A(_0246_),
    .B1(_0212_),
    .B2(_0211_),
    .ZN(_0247_));
 INV_X1 _3922_ (.A(_0186_),
    .ZN(_0248_));
 NAND2_X1 _3923_ (.A1(_0248_),
    .A2(_0208_),
    .ZN(_0249_));
 OAI21_X1 _3924_ (.A(_0249_),
    .B1(_0210_),
    .B2(_0184_),
    .ZN(_0250_));
 NAND2_X1 _3925_ (.A1(_0158_),
    .A2(_0209_),
    .ZN(_0251_));
 AOI21_X1 _3926_ (.A(_0251_),
    .B1(_2850_),
    .B2(_2953_),
    .ZN(_0252_));
 NAND4_X1 _3927_ (.A1(_2757_),
    .A2(_2846_),
    .A3(_0158_),
    .A4(_0209_),
    .ZN(_0253_));
 NAND3_X1 _3928_ (.A1(_2553_),
    .A2(_2614_),
    .A3(_2681_),
    .ZN(_0254_));
 AOI21_X1 _3929_ (.A(_0253_),
    .B1(_0254_),
    .B2(_2700_),
    .ZN(_0255_));
 NOR2_X1 _3930_ (.A1(_2485_),
    .A2(_2544_),
    .ZN(_0256_));
 NAND3_X1 _3931_ (.A1(_0256_),
    .A2(_2614_),
    .A3(_2681_),
    .ZN(_0257_));
 NOR3_X1 _3932_ (.A1(_2425_),
    .A2(_0257_),
    .A3(_0253_),
    .ZN(_0258_));
 NOR4_X1 _3933_ (.A1(_0250_),
    .A2(_0252_),
    .A3(_0255_),
    .A4(_0258_),
    .ZN(_0259_));
 NAND3_X1 _3934_ (.A1(\section_2.xn2[10] ),
    .A2(\section_2.xn2[9] ),
    .A3(_0207_),
    .ZN(_0260_));
 OAI21_X1 _3935_ (.A(_0260_),
    .B1(_0206_),
    .B2(_0189_),
    .ZN(_0261_));
 NOR2_X1 _3936_ (.A1(_0031_),
    .A2(_0152_),
    .ZN(_0262_));
 NAND2_X1 _3937_ (.A1(_0262_),
    .A2(_0205_),
    .ZN(_0263_));
 NOR2_X1 _3938_ (.A1(_0031_),
    .A2(_0205_),
    .ZN(_0264_));
 NAND2_X1 _3939_ (.A1(_0148_),
    .A2(_0201_),
    .ZN(_0265_));
 INV_X1 _3940_ (.A(_0204_),
    .ZN(_0266_));
 OAI21_X1 _3941_ (.A(_0265_),
    .B1(_0202_),
    .B2(_0266_),
    .ZN(_0267_));
 INV_X1 _3942_ (.A(_0192_),
    .ZN(_0268_));
 NAND2_X1 _3943_ (.A1(_0268_),
    .A2(_0200_),
    .ZN(_0269_));
 AOI21_X1 _3944_ (.A(_2717_),
    .B1(_0195_),
    .B2(_0197_),
    .ZN(_0270_));
 AOI21_X1 _3945_ (.A(_0198_),
    .B1(_0143_),
    .B2(\section_1.yn2[10] ),
    .ZN(_0271_));
 OR2_X1 _3946_ (.A1(_0270_),
    .A2(_0271_),
    .ZN(_0272_));
 INV_X1 _3947_ (.A(_0272_),
    .ZN(_0273_));
 NOR2_X1 _3948_ (.A1(_2717_),
    .A2(_0198_),
    .ZN(_0274_));
 XNOR2_X1 _3949_ (.A(\coll_reg[10] ),
    .B(_0004_),
    .ZN(_0275_));
 XNOR2_X1 _3950_ (.A(_0274_),
    .B(_0275_),
    .ZN(_0276_));
 XNOR2_X1 _3951_ (.A(_0273_),
    .B(_0276_),
    .ZN(_0277_));
 XOR2_X1 _3952_ (.A(_0269_),
    .B(_0277_),
    .Z(_0278_));
 XNOR2_X1 _3953_ (.A(_0267_),
    .B(_0278_),
    .ZN(_0279_));
 XNOR2_X1 _3954_ (.A(_2639_),
    .B(_0279_),
    .ZN(_0280_));
 XNOR2_X1 _3955_ (.A(_0264_),
    .B(_0280_),
    .ZN(_0281_));
 XNOR2_X1 _3956_ (.A(_0263_),
    .B(_0281_),
    .ZN(_0282_));
 XNOR2_X1 _3957_ (.A(\section_2.xn2[10] ),
    .B(_0282_),
    .ZN(_0283_));
 XNOR2_X1 _3958_ (.A(_0261_),
    .B(_0283_),
    .ZN(_0284_));
 XNOR2_X1 _3959_ (.A(_0259_),
    .B(_0284_),
    .ZN(_0285_));
 XOR2_X1 _3960_ (.A(_0247_),
    .B(_0285_),
    .Z(_0286_));
 XOR2_X1 _3961_ (.A(_0245_),
    .B(_0286_),
    .Z(_0287_));
 XNOR2_X1 _3962_ (.A(_0239_),
    .B(_0287_),
    .ZN(_0288_));
 XNOR2_X1 _3963_ (.A(_0237_),
    .B(_0288_),
    .ZN(_0289_));
 XOR2_X1 _3964_ (.A(_0236_),
    .B(_0289_),
    .Z(_0290_));
 XOR2_X1 _3965_ (.A(_0234_),
    .B(_0290_),
    .Z(_0291_));
 XNOR2_X1 _3966_ (.A(_0169_),
    .B(_0291_),
    .ZN(_0292_));
 XNOR2_X1 _3967_ (.A(_0233_),
    .B(_0292_),
    .ZN(_0293_));
 XNOR2_X1 _3968_ (.A(_0229_),
    .B(_0293_),
    .ZN(_0294_));
 XNOR2_X1 _3969_ (.A(_0231_),
    .B(_0294_),
    .ZN(_0295_));
 NOR2_X1 _3970_ (.A1(_0230_),
    .A2(_0295_),
    .ZN(_0296_));
 INV_X1 _3971_ (.A(\section_2.yn2[6] ),
    .ZN(_0297_));
 NAND2_X1 _3972_ (.A1(\section_2.yn2[10] ),
    .A2(\section_2.yn2[8] ),
    .ZN(_0298_));
 XNOR2_X1 _3973_ (.A(_0297_),
    .B(_0298_),
    .ZN(_0299_));
 XOR2_X1 _3974_ (.A(_0230_),
    .B(_0295_),
    .Z(_0300_));
 AOI21_X1 _3975_ (.A(_0296_),
    .B1(_0299_),
    .B2(_0300_),
    .ZN(_0301_));
 NAND2_X1 _3976_ (.A1(\section_2.yn2[10] ),
    .A2(\section_2.yn2[9] ),
    .ZN(_0302_));
 XOR2_X1 _3977_ (.A(\section_2.yn2[7] ),
    .B(_0302_),
    .Z(_0303_));
 INV_X1 _3978_ (.A(_0002_),
    .ZN(_0304_));
 AND3_X1 _3979_ (.A1(_0304_),
    .A2(_0227_),
    .A3(_0293_),
    .ZN(_0305_));
 AOI21_X1 _3980_ (.A(_0305_),
    .B1(_0294_),
    .B2(_0231_),
    .ZN(_0306_));
 NAND2_X1 _3981_ (.A1(_0304_),
    .A2(_0293_),
    .ZN(_0307_));
 INV_X1 _3982_ (.A(_0236_),
    .ZN(_0308_));
 NAND2_X1 _3983_ (.A1(_0308_),
    .A2(_0289_),
    .ZN(_0309_));
 AND2_X1 _3984_ (.A1(_0239_),
    .A2(_0287_),
    .ZN(_0310_));
 NOR3_X1 _3985_ (.A1(z[6]),
    .A2(_2947_),
    .A3(_0288_),
    .ZN(_0311_));
 AND3_X1 _3986_ (.A1(z[10]),
    .A2(_0161_),
    .A3(_0213_),
    .ZN(_0312_));
 AOI22_X1 _3987_ (.A1(_0312_),
    .A2(_0285_),
    .B1(_0286_),
    .B2(_0245_),
    .ZN(_0313_));
 NOR2_X1 _3988_ (.A1(z[8]),
    .A2(_0243_),
    .ZN(_0314_));
 OR2_X1 _3989_ (.A1(z[8]),
    .A2(z[7]),
    .ZN(_0315_));
 NAND2_X1 _3990_ (.A1(z[8]),
    .A2(z[7]),
    .ZN(_0316_));
 AOI22_X1 _3991_ (.A1(z[7]),
    .A2(z[6]),
    .B1(_0315_),
    .B2(_0316_),
    .ZN(_0317_));
 NOR2_X1 _3992_ (.A1(_0314_),
    .A2(_0317_),
    .ZN(_0318_));
 OAI211_X1 _3993_ (.A(z[10]),
    .B(_0285_),
    .C1(_0212_),
    .C2(_0211_),
    .ZN(_0319_));
 NAND2_X1 _3994_ (.A1(_0261_),
    .A2(_0283_),
    .ZN(_0320_));
 OAI21_X1 _3995_ (.A(_0320_),
    .B1(_0284_),
    .B2(_0259_),
    .ZN(_0321_));
 NOR2_X1 _3996_ (.A1(_0263_),
    .A2(_0281_),
    .ZN(_0322_));
 NAND2_X1 _3997_ (.A1(_0263_),
    .A2(_0281_),
    .ZN(_0323_));
 AOI21_X1 _3998_ (.A(_0322_),
    .B1(_0323_),
    .B2(\section_2.xn2[10] ),
    .ZN(_0324_));
 NAND2_X1 _3999_ (.A1(_0279_),
    .A2(_0264_),
    .ZN(_0325_));
 NOR2_X1 _4000_ (.A1(_0031_),
    .A2(_0279_),
    .ZN(_0326_));
 NOR2_X1 _4001_ (.A1(_0269_),
    .A2(_0277_),
    .ZN(_0327_));
 AOI21_X1 _4002_ (.A(_0327_),
    .B1(_0278_),
    .B2(_0267_),
    .ZN(_0328_));
 NAND2_X1 _4003_ (.A1(_0273_),
    .A2(_0276_),
    .ZN(_0329_));
 INV_X1 _4004_ (.A(net89),
    .ZN(_0330_));
 MUX2_X1 _4005_ (.A(_2717_),
    .B(_0270_),
    .S(_0330_),
    .Z(_0331_));
 NOR2_X1 _4006_ (.A1(\section_1.yn2[10] ),
    .A2(\coll_reg[10] ),
    .ZN(_0332_));
 XNOR2_X1 _4007_ (.A(_0004_),
    .B(_0332_),
    .ZN(_0333_));
 XOR2_X1 _4008_ (.A(_0331_),
    .B(_0333_),
    .Z(_0334_));
 XNOR2_X1 _4009_ (.A(_0329_),
    .B(_0334_),
    .ZN(_0335_));
 XNOR2_X1 _4010_ (.A(_0328_),
    .B(_0335_),
    .ZN(_0336_));
 XNOR2_X1 _4011_ (.A(_0031_),
    .B(_0336_),
    .ZN(_0337_));
 XNOR2_X1 _4012_ (.A(_0326_),
    .B(_0337_),
    .ZN(_0338_));
 XOR2_X1 _4013_ (.A(_0325_),
    .B(_0338_),
    .Z(_0339_));
 XNOR2_X1 _4014_ (.A(\section_2.xn2[10] ),
    .B(_0339_),
    .ZN(_0340_));
 XOR2_X1 _4015_ (.A(_0324_),
    .B(_0340_),
    .Z(_0341_));
 XNOR2_X1 _4016_ (.A(_0321_),
    .B(_0341_),
    .ZN(_0342_));
 XOR2_X1 _4017_ (.A(_0319_),
    .B(_0342_),
    .Z(_0343_));
 XOR2_X1 _4018_ (.A(_0318_),
    .B(_0343_),
    .Z(_0344_));
 XNOR2_X1 _4019_ (.A(_0313_),
    .B(_0344_),
    .ZN(_0345_));
 XOR2_X1 _4020_ (.A(_0241_),
    .B(_0345_),
    .Z(_0346_));
 OR3_X1 _4021_ (.A1(_0310_),
    .A2(_0311_),
    .A3(_0346_),
    .ZN(_0347_));
 OAI21_X1 _4022_ (.A(_0346_),
    .B1(_0311_),
    .B2(_0310_),
    .ZN(_0348_));
 NAND2_X1 _4023_ (.A1(_0347_),
    .A2(_0348_),
    .ZN(_0349_));
 XOR2_X1 _4024_ (.A(_0309_),
    .B(_0349_),
    .Z(_0350_));
 NAND2_X1 _4025_ (.A1(_0219_),
    .A2(_0291_),
    .ZN(_0351_));
 AOI21_X1 _4026_ (.A(_0351_),
    .B1(_0224_),
    .B2(_0223_),
    .ZN(_0352_));
 NOR2_X1 _4027_ (.A1(_0234_),
    .A2(_0290_),
    .ZN(_0353_));
 AOI21_X1 _4028_ (.A(_0353_),
    .B1(_0291_),
    .B2(_0232_),
    .ZN(_0354_));
 INV_X1 _4029_ (.A(_0354_),
    .ZN(_0355_));
 OR2_X1 _4030_ (.A1(_0352_),
    .A2(_0355_),
    .ZN(_0356_));
 XOR2_X1 _4031_ (.A(_0350_),
    .B(_0356_),
    .Z(_0357_));
 XNOR2_X1 _4032_ (.A(_0169_),
    .B(_0357_),
    .ZN(_0358_));
 XNOR2_X1 _4033_ (.A(_0307_),
    .B(_0358_),
    .ZN(_0359_));
 XOR2_X1 _4034_ (.A(_0306_),
    .B(_0359_),
    .Z(_0360_));
 XNOR2_X1 _4035_ (.A(_0303_),
    .B(_0360_),
    .ZN(_0361_));
 NOR2_X1 _4036_ (.A1(_0301_),
    .A2(_0361_),
    .ZN(_0362_));
 XOR2_X1 _4037_ (.A(_0301_),
    .B(_0361_),
    .Z(_0363_));
 NOR2_X1 _4038_ (.A1(\section_2.yn2[6] ),
    .A2(_0298_),
    .ZN(_0364_));
 AOI21_X1 _4039_ (.A(_0362_),
    .B1(_0363_),
    .B2(_0364_),
    .ZN(_0365_));
 OR2_X1 _4040_ (.A1(\section_2.yn2[7] ),
    .A2(_0302_),
    .ZN(_0366_));
 NOR2_X1 _4041_ (.A1(_0306_),
    .A2(_0359_),
    .ZN(_0367_));
 AOI21_X1 _4042_ (.A(_0367_),
    .B1(_0360_),
    .B2(_0303_),
    .ZN(_0368_));
 NAND2_X1 _4043_ (.A1(_0304_),
    .A2(_0358_),
    .ZN(_0369_));
 NOR2_X1 _4044_ (.A1(_0293_),
    .A2(_0369_),
    .ZN(_0370_));
 NOR2_X1 _4045_ (.A1(_0309_),
    .A2(_0349_),
    .ZN(_0371_));
 INV_X1 _4046_ (.A(_0371_),
    .ZN(_0372_));
 OAI21_X1 _4047_ (.A(_0350_),
    .B1(_0352_),
    .B2(_0355_),
    .ZN(_0373_));
 INV_X1 _4048_ (.A(_0313_),
    .ZN(_0374_));
 NAND2_X1 _4049_ (.A1(_0374_),
    .A2(_0344_),
    .ZN(_0375_));
 NAND2_X1 _4050_ (.A1(_0241_),
    .A2(_0345_),
    .ZN(_0376_));
 NAND2_X1 _4051_ (.A1(_0375_),
    .A2(_0376_),
    .ZN(_0377_));
 NAND3_X1 _4052_ (.A1(z[10]),
    .A2(_0285_),
    .A3(_0342_),
    .ZN(_0378_));
 NOR2_X1 _4053_ (.A1(_0213_),
    .A2(_0378_),
    .ZN(_0379_));
 AOI21_X1 _4054_ (.A(_0379_),
    .B1(_0343_),
    .B2(_0318_),
    .ZN(_0380_));
 XOR2_X1 _4055_ (.A(z[9]),
    .B(z[8]),
    .Z(_0381_));
 XNOR2_X1 _4056_ (.A(_0316_),
    .B(_0381_),
    .ZN(_0382_));
 NOR2_X1 _4057_ (.A1(_0324_),
    .A2(_0340_),
    .ZN(_0383_));
 AOI21_X1 _4058_ (.A(_0383_),
    .B1(_0341_),
    .B2(_0321_),
    .ZN(_0384_));
 NOR2_X1 _4059_ (.A1(_0325_),
    .A2(_0336_),
    .ZN(_0385_));
 AOI21_X1 _4060_ (.A(_0385_),
    .B1(_0339_),
    .B2(\section_2.xn2[10] ),
    .ZN(_0386_));
 INV_X1 _4061_ (.A(_0335_),
    .ZN(_0387_));
 XNOR2_X1 _4062_ (.A(_0328_),
    .B(_0387_),
    .ZN(_0388_));
 NAND2_X1 _4063_ (.A1(_0326_),
    .A2(_0388_),
    .ZN(_0389_));
 NAND3_X1 _4064_ (.A1(_0273_),
    .A2(_0276_),
    .A3(_0334_),
    .ZN(_0390_));
 NOR3_X1 _4065_ (.A1(_2717_),
    .A2(_0330_),
    .A3(_0144_),
    .ZN(_0391_));
 AOI21_X1 _4066_ (.A(_0391_),
    .B1(_0333_),
    .B2(_0331_),
    .ZN(_0392_));
 OAI211_X1 _4067_ (.A(_0390_),
    .B(_0392_),
    .C1(_0387_),
    .C2(_0328_),
    .ZN(_0393_));
 XOR2_X1 _4068_ (.A(\section_2.xn2[10] ),
    .B(_0393_),
    .Z(_0394_));
 OR2_X1 _4069_ (.A1(_0389_),
    .A2(_0394_),
    .ZN(_0395_));
 NOR2_X1 _4070_ (.A1(_0031_),
    .A2(_0388_),
    .ZN(_0396_));
 XOR2_X1 _4071_ (.A(_0396_),
    .B(_0394_),
    .Z(_0397_));
 NAND2_X1 _4072_ (.A1(_0389_),
    .A2(_0397_),
    .ZN(_0398_));
 NAND2_X1 _4073_ (.A1(_0395_),
    .A2(_0398_),
    .ZN(_0399_));
 XOR2_X1 _4074_ (.A(\section_2.xn2[10] ),
    .B(_0399_),
    .Z(_0400_));
 XNOR2_X1 _4075_ (.A(_0386_),
    .B(_0400_),
    .ZN(_0401_));
 XNOR2_X1 _4076_ (.A(_0384_),
    .B(_0401_),
    .ZN(_0402_));
 XOR2_X1 _4077_ (.A(_0378_),
    .B(_0402_),
    .Z(_0403_));
 XOR2_X1 _4078_ (.A(_0382_),
    .B(_0403_),
    .Z(_0404_));
 XOR2_X1 _4079_ (.A(_0380_),
    .B(_0404_),
    .Z(_0405_));
 XNOR2_X1 _4080_ (.A(_0314_),
    .B(_0405_),
    .ZN(_0406_));
 XNOR2_X1 _4081_ (.A(_0377_),
    .B(_0406_),
    .ZN(_0407_));
 XOR2_X1 _4082_ (.A(_0348_),
    .B(_0407_),
    .Z(_0408_));
 INV_X1 _4083_ (.A(_0408_),
    .ZN(_0409_));
 AND3_X1 _4084_ (.A1(_0372_),
    .A2(_0373_),
    .A3(_0409_),
    .ZN(_0410_));
 AOI21_X1 _4085_ (.A(_0409_),
    .B1(_0373_),
    .B2(_0372_),
    .ZN(_0411_));
 OR2_X1 _4086_ (.A1(_0410_),
    .A2(_0411_),
    .ZN(_0412_));
 XNOR2_X1 _4087_ (.A(_0169_),
    .B(_0412_),
    .ZN(_0413_));
 XNOR2_X1 _4088_ (.A(_0369_),
    .B(_0413_),
    .ZN(_0414_));
 XNOR2_X1 _4089_ (.A(_0370_),
    .B(_0414_),
    .ZN(_0415_));
 XNOR2_X1 _4090_ (.A(_1264_),
    .B(_0415_),
    .ZN(_0416_));
 XNOR2_X1 _4091_ (.A(_0368_),
    .B(_0416_),
    .ZN(_0417_));
 XNOR2_X1 _4092_ (.A(_0366_),
    .B(_0417_),
    .ZN(_0418_));
 NOR2_X1 _4093_ (.A1(_0365_),
    .A2(_0418_),
    .ZN(_0419_));
 XNOR2_X1 _4094_ (.A(_2861_),
    .B(_2934_),
    .ZN(_0420_));
 XNOR2_X1 _4095_ (.A(_0169_),
    .B(_0420_),
    .ZN(_0421_));
 NOR2_X1 _4096_ (.A1(_0002_),
    .A2(_0421_),
    .ZN(_0422_));
 XOR2_X1 _4097_ (.A(_0171_),
    .B(_0422_),
    .Z(_0423_));
 INV_X1 _4098_ (.A(_0423_),
    .ZN(_0424_));
 XOR2_X1 _4099_ (.A(\section_2.yn2[10] ),
    .B(\section_2.yn2[7] ),
    .Z(_0425_));
 AOI22_X1 _4100_ (.A1(_0173_),
    .A2(_0421_),
    .B1(_0424_),
    .B2(_0425_),
    .ZN(_0426_));
 XNOR2_X1 _4101_ (.A(_1264_),
    .B(_0228_),
    .ZN(_0427_));
 NOR2_X1 _4102_ (.A1(_0426_),
    .A2(_0427_),
    .ZN(_0428_));
 INV_X1 _4103_ (.A(\section_2.yn2[5] ),
    .ZN(_0429_));
 NAND2_X1 _4104_ (.A1(\section_2.yn2[10] ),
    .A2(\section_2.yn2[7] ),
    .ZN(_0430_));
 XNOR2_X1 _4105_ (.A(_0429_),
    .B(_0430_),
    .ZN(_0431_));
 XOR2_X1 _4106_ (.A(_0426_),
    .B(_0427_),
    .Z(_0432_));
 AOI21_X1 _4107_ (.A(_0428_),
    .B1(_0431_),
    .B2(_0432_),
    .ZN(_0433_));
 XNOR2_X1 _4108_ (.A(_0299_),
    .B(_0300_),
    .ZN(_0434_));
 NOR2_X1 _4109_ (.A1(_0433_),
    .A2(_0434_),
    .ZN(_0435_));
 XOR2_X1 _4110_ (.A(_0433_),
    .B(_0434_),
    .Z(_0436_));
 NOR2_X1 _4111_ (.A1(\section_2.yn2[5] ),
    .A2(_0430_),
    .ZN(_0437_));
 AOI21_X1 _4112_ (.A(_0435_),
    .B1(_0436_),
    .B2(_0437_),
    .ZN(_0438_));
 XNOR2_X1 _4113_ (.A(_0364_),
    .B(_0363_),
    .ZN(_0439_));
 NOR2_X1 _4114_ (.A1(_0438_),
    .A2(_0439_),
    .ZN(_0440_));
 XOR2_X1 _4115_ (.A(_0438_),
    .B(_0439_),
    .Z(_0441_));
 INV_X1 _4116_ (.A(\section_2.yn2[10] ),
    .ZN(_0442_));
 XNOR2_X1 _4117_ (.A(_0442_),
    .B(_0420_),
    .ZN(_0443_));
 AND2_X1 _4118_ (.A1(_2872_),
    .A2(_2873_),
    .ZN(_0444_));
 OAI21_X1 _4119_ (.A(_2876_),
    .B1(_2877_),
    .B2(_2878_),
    .ZN(_0445_));
 AOI21_X1 _4120_ (.A(_0444_),
    .B1(_0445_),
    .B2(_2794_),
    .ZN(_0446_));
 OAI221_X1 _4121_ (.A(_2894_),
    .B1(_2931_),
    .B2(_2932_),
    .C1(_2881_),
    .C2(_0446_),
    .ZN(_0447_));
 NAND3_X1 _4122_ (.A1(_2794_),
    .A2(_0444_),
    .A3(_0445_),
    .ZN(_0448_));
 NAND3_X1 _4123_ (.A1(_2880_),
    .A2(_0448_),
    .A3(_2933_),
    .ZN(_0449_));
 NAND3_X1 _4124_ (.A1(_0304_),
    .A2(_0447_),
    .A3(_0449_),
    .ZN(_0450_));
 AOI21_X1 _4125_ (.A(_2933_),
    .B1(_0448_),
    .B2(_2880_),
    .ZN(_0451_));
 AND3_X1 _4126_ (.A1(_2880_),
    .A2(_0448_),
    .A3(_2933_),
    .ZN(_0452_));
 OAI21_X1 _4127_ (.A(_0002_),
    .B1(_0451_),
    .B2(_0452_),
    .ZN(_0453_));
 NAND3_X1 _4128_ (.A1(_0231_),
    .A2(_0450_),
    .A3(_0453_),
    .ZN(_0454_));
 AOI21_X1 _4129_ (.A(_0443_),
    .B1(_0450_),
    .B2(_0454_),
    .ZN(_0455_));
 XOR2_X1 _4130_ (.A(_0026_),
    .B(_0302_),
    .Z(_0456_));
 AOI21_X1 _4131_ (.A(_0304_),
    .B1(_0447_),
    .B2(_0449_),
    .ZN(_0457_));
 INV_X1 _4132_ (.A(_0231_),
    .ZN(_0458_));
 OAI21_X1 _4133_ (.A(_0450_),
    .B1(_0457_),
    .B2(_0458_),
    .ZN(_0459_));
 XNOR2_X1 _4134_ (.A(_0443_),
    .B(_0459_),
    .ZN(_0460_));
 AOI21_X1 _4135_ (.A(_0455_),
    .B1(_0456_),
    .B2(_0460_),
    .ZN(_0461_));
 XOR2_X1 _4136_ (.A(_0425_),
    .B(_0423_),
    .Z(_0462_));
 NOR2_X1 _4137_ (.A1(_0461_),
    .A2(_0462_),
    .ZN(_0463_));
 NOR2_X1 _4138_ (.A1(_0026_),
    .A2(_0302_),
    .ZN(_0464_));
 XNOR2_X1 _4139_ (.A(\section_2.yn2[4] ),
    .B(_0464_),
    .ZN(_0465_));
 XOR2_X1 _4140_ (.A(_0461_),
    .B(_0462_),
    .Z(_0466_));
 AOI21_X1 _4141_ (.A(_0463_),
    .B1(_0465_),
    .B2(_0466_),
    .ZN(_0467_));
 XNOR2_X1 _4142_ (.A(_0431_),
    .B(_0432_),
    .ZN(_0468_));
 NOR2_X1 _4143_ (.A1(_0467_),
    .A2(_0468_),
    .ZN(_0469_));
 XOR2_X1 _4144_ (.A(_0467_),
    .B(_0468_),
    .Z(_0470_));
 NOR3_X1 _4145_ (.A1(\section_2.yn2[4] ),
    .A2(_0026_),
    .A3(_0302_),
    .ZN(_0471_));
 AOI21_X1 _4146_ (.A(_0469_),
    .B1(_0470_),
    .B2(_0471_),
    .ZN(_0472_));
 XNOR2_X1 _4147_ (.A(_0437_),
    .B(_0436_),
    .ZN(_0473_));
 NOR2_X1 _4148_ (.A1(_0472_),
    .A2(_0473_),
    .ZN(_0474_));
 AOI21_X1 _4149_ (.A(_0440_),
    .B1(_0441_),
    .B2(_0474_),
    .ZN(_0475_));
 XOR2_X1 _4150_ (.A(_0472_),
    .B(_0473_),
    .Z(_0476_));
 NAND2_X1 _4151_ (.A1(_0441_),
    .A2(_0476_),
    .ZN(_0477_));
 XNOR2_X1 _4152_ (.A(_0456_),
    .B(_0460_),
    .ZN(_0478_));
 NOR3_X1 _4153_ (.A1(_0002_),
    .A2(_0451_),
    .A3(_0452_),
    .ZN(_0479_));
 NOR3_X1 _4154_ (.A1(_0458_),
    .A2(_0479_),
    .A3(_0457_),
    .ZN(_0480_));
 XOR2_X1 _4155_ (.A(_2904_),
    .B(_2930_),
    .Z(_0481_));
 OR2_X1 _4156_ (.A1(\section_2.yn2[10] ),
    .A2(_0481_),
    .ZN(_0482_));
 XNOR2_X1 _4157_ (.A(_2931_),
    .B(_2932_),
    .ZN(_0483_));
 XNOR2_X1 _4158_ (.A(_0169_),
    .B(_0483_),
    .ZN(_0484_));
 AND2_X1 _4159_ (.A1(_0482_),
    .A2(_0484_),
    .ZN(_0485_));
 XOR2_X1 _4160_ (.A(\section_2.yn2[9] ),
    .B(\section_2.yn2[8] ),
    .Z(_0486_));
 OR2_X1 _4161_ (.A1(_0482_),
    .A2(_0484_),
    .ZN(_0487_));
 AOI21_X1 _4162_ (.A(_0485_),
    .B1(_0486_),
    .B2(_0487_),
    .ZN(_0488_));
 AOI21_X1 _4163_ (.A(_0231_),
    .B1(_0450_),
    .B2(_0453_),
    .ZN(_0489_));
 OR3_X1 _4164_ (.A1(_0480_),
    .A2(_0488_),
    .A3(_0489_),
    .ZN(_0490_));
 INV_X1 _4165_ (.A(_0028_),
    .ZN(_0491_));
 NAND2_X1 _4166_ (.A1(\section_2.yn2[9] ),
    .A2(\section_2.yn2[8] ),
    .ZN(_0492_));
 XNOR2_X1 _4167_ (.A(_0491_),
    .B(_0492_),
    .ZN(_0493_));
 OAI21_X1 _4168_ (.A(_0488_),
    .B1(_0489_),
    .B2(_0480_),
    .ZN(_0494_));
 NAND3_X1 _4169_ (.A1(_0490_),
    .A2(_0493_),
    .A3(_0494_),
    .ZN(_0495_));
 AOI21_X1 _4170_ (.A(_0478_),
    .B1(_0495_),
    .B2(_0490_),
    .ZN(_0496_));
 NOR3_X1 _4171_ (.A1(\section_2.yn2[3] ),
    .A2(_0028_),
    .A3(_0492_),
    .ZN(_0497_));
 INV_X1 _4172_ (.A(\section_2.yn2[3] ),
    .ZN(_0498_));
 INV_X1 _4173_ (.A(_0492_),
    .ZN(_0499_));
 AOI21_X1 _4174_ (.A(_0498_),
    .B1(_0491_),
    .B2(_0499_),
    .ZN(_0500_));
 NOR2_X1 _4175_ (.A1(_0497_),
    .A2(_0500_),
    .ZN(_0501_));
 INV_X1 _4176_ (.A(_0493_),
    .ZN(_0502_));
 OAI21_X1 _4177_ (.A(_0458_),
    .B1(_0479_),
    .B2(_0457_),
    .ZN(_0503_));
 AOI221_X1 _4178_ (.A(_0485_),
    .B1(_0486_),
    .B2(_0487_),
    .C1(_0503_),
    .C2(_0454_),
    .ZN(_0504_));
 OAI21_X1 _4179_ (.A(_0490_),
    .B1(_0502_),
    .B2(_0504_),
    .ZN(_0505_));
 XNOR2_X1 _4180_ (.A(_0505_),
    .B(_0478_),
    .ZN(_0506_));
 AOI21_X1 _4181_ (.A(_0496_),
    .B1(_0501_),
    .B2(_0506_),
    .ZN(_0507_));
 XNOR2_X1 _4182_ (.A(_0465_),
    .B(_0466_),
    .ZN(_0508_));
 NOR2_X1 _4183_ (.A1(_0507_),
    .A2(_0508_),
    .ZN(_0509_));
 XOR2_X1 _4184_ (.A(_0507_),
    .B(_0508_),
    .Z(_0510_));
 AOI21_X1 _4185_ (.A(_0509_),
    .B1(_0510_),
    .B2(_0497_),
    .ZN(_0511_));
 XNOR2_X1 _4186_ (.A(_0471_),
    .B(_0470_),
    .ZN(_0512_));
 NOR2_X1 _4187_ (.A1(_0511_),
    .A2(_0512_),
    .ZN(_0513_));
 XOR2_X1 _4188_ (.A(_0511_),
    .B(_0512_),
    .Z(_0514_));
 XOR2_X1 _4189_ (.A(_0497_),
    .B(_0510_),
    .Z(_0515_));
 INV_X1 _4190_ (.A(\section_2.yn2[4] ),
    .ZN(_0516_));
 AOI21_X1 _4191_ (.A(_0499_),
    .B1(_0486_),
    .B2(\section_2.yn2[7] ),
    .ZN(_0517_));
 OR2_X1 _4192_ (.A1(_0516_),
    .A2(_0517_),
    .ZN(_0518_));
 NOR2_X1 _4193_ (.A1(\section_2.yn2[2] ),
    .A2(_0518_),
    .ZN(_0519_));
 NOR3_X1 _4194_ (.A1(_0480_),
    .A2(_0488_),
    .A3(_0489_),
    .ZN(_0520_));
 NOR3_X1 _4195_ (.A1(_0520_),
    .A2(_0502_),
    .A3(_0504_),
    .ZN(_0521_));
 XOR2_X1 _4196_ (.A(_2928_),
    .B(_2929_),
    .Z(_0522_));
 NAND2_X1 _4197_ (.A1(\section_2.yn2[9] ),
    .A2(_0522_),
    .ZN(_0523_));
 XNOR2_X1 _4198_ (.A(\section_2.yn2[9] ),
    .B(_0522_),
    .ZN(_0524_));
 INV_X1 _4199_ (.A(\section_2.yn2[8] ),
    .ZN(_0525_));
 OAI21_X1 _4200_ (.A(_0523_),
    .B1(_0524_),
    .B2(_0525_),
    .ZN(_0526_));
 XNOR2_X1 _4201_ (.A(_0304_),
    .B(_0481_),
    .ZN(_0527_));
 NAND2_X1 _4202_ (.A1(_0526_),
    .A2(_0527_),
    .ZN(_0528_));
 XNOR2_X1 _4203_ (.A(\section_2.yn2[7] ),
    .B(_0486_),
    .ZN(_0529_));
 XNOR2_X1 _4204_ (.A(_0526_),
    .B(_0527_),
    .ZN(_0530_));
 OAI21_X1 _4205_ (.A(_0528_),
    .B1(_0529_),
    .B2(_0530_),
    .ZN(_0531_));
 XNOR2_X1 _4206_ (.A(_0482_),
    .B(_0484_),
    .ZN(_0532_));
 XNOR2_X1 _4207_ (.A(_0486_),
    .B(_0532_),
    .ZN(_0533_));
 AND2_X1 _4208_ (.A1(_0531_),
    .A2(_0533_),
    .ZN(_0534_));
 XNOR2_X1 _4209_ (.A(\section_2.yn2[4] ),
    .B(_0517_),
    .ZN(_0535_));
 OR2_X1 _4210_ (.A1(_0531_),
    .A2(_0533_),
    .ZN(_0536_));
 AOI21_X1 _4211_ (.A(_0534_),
    .B1(_0535_),
    .B2(_0536_),
    .ZN(_0537_));
 AOI21_X1 _4212_ (.A(_0493_),
    .B1(_0494_),
    .B2(_0490_),
    .ZN(_0538_));
 NOR3_X1 _4213_ (.A1(_0521_),
    .A2(_0537_),
    .A3(_0538_),
    .ZN(_0539_));
 INV_X1 _4214_ (.A(\section_2.yn2[2] ),
    .ZN(_0540_));
 XNOR2_X1 _4215_ (.A(_0540_),
    .B(_0518_),
    .ZN(_0541_));
 OAI21_X1 _4216_ (.A(_0537_),
    .B1(_0538_),
    .B2(_0521_),
    .ZN(_0542_));
 AOI21_X1 _4217_ (.A(_0539_),
    .B1(_0541_),
    .B2(_0542_),
    .ZN(_0543_));
 XNOR2_X1 _4218_ (.A(_0501_),
    .B(_0506_),
    .ZN(_0544_));
 XOR2_X1 _4219_ (.A(_0543_),
    .B(_0544_),
    .Z(_0545_));
 AND2_X1 _4220_ (.A1(_0519_),
    .A2(_0545_),
    .ZN(_0546_));
 NOR2_X1 _4221_ (.A1(_0543_),
    .A2(_0544_),
    .ZN(_0547_));
 OAI21_X1 _4222_ (.A(_0515_),
    .B1(_0546_),
    .B2(_0547_),
    .ZN(_0548_));
 OR3_X1 _4223_ (.A1(_0547_),
    .A2(_0546_),
    .A3(_0515_),
    .ZN(_0549_));
 NAND2_X1 _4224_ (.A1(_0548_),
    .A2(_0549_),
    .ZN(_0550_));
 INV_X1 _4225_ (.A(_0541_),
    .ZN(_0551_));
 OAI21_X1 _4226_ (.A(_0502_),
    .B1(_0504_),
    .B2(_0520_),
    .ZN(_0552_));
 AOI221_X1 _4227_ (.A(_0534_),
    .B1(_0535_),
    .B2(_0536_),
    .C1(_0552_),
    .C2(_0495_),
    .ZN(_0553_));
 NOR3_X1 _4228_ (.A1(_0539_),
    .A2(_0551_),
    .A3(_0553_),
    .ZN(_0554_));
 XNOR2_X1 _4229_ (.A(_0531_),
    .B(_0533_),
    .ZN(_0555_));
 XOR2_X1 _4230_ (.A(_0535_),
    .B(_0555_),
    .Z(_0556_));
 XNOR2_X1 _4231_ (.A(_0525_),
    .B(_0524_),
    .ZN(_0557_));
 OAI21_X1 _4232_ (.A(_2914_),
    .B1(_2926_),
    .B2(_2927_),
    .ZN(_0558_));
 XOR2_X1 _4233_ (.A(_2916_),
    .B(_0558_),
    .Z(_0559_));
 XNOR2_X1 _4234_ (.A(_0525_),
    .B(_0559_),
    .ZN(_0560_));
 INV_X1 _4235_ (.A(_0560_),
    .ZN(_0561_));
 NAND2_X1 _4236_ (.A1(\section_2.yn2[7] ),
    .A2(_0561_),
    .ZN(_0562_));
 OR2_X1 _4237_ (.A1(_0525_),
    .A2(_0559_),
    .ZN(_0563_));
 AOI21_X1 _4238_ (.A(_0557_),
    .B1(_0562_),
    .B2(_0563_),
    .ZN(_0564_));
 XOR2_X1 _4239_ (.A(\section_2.yn2[7] ),
    .B(\section_2.yn2[6] ),
    .Z(_0565_));
 NAND3_X1 _4240_ (.A1(_0563_),
    .A2(_0562_),
    .A3(_0557_),
    .ZN(_0566_));
 AOI21_X1 _4241_ (.A(_0564_),
    .B1(_0565_),
    .B2(_0566_),
    .ZN(_0567_));
 XOR2_X1 _4242_ (.A(_0529_),
    .B(_0530_),
    .Z(_0568_));
 XNOR2_X1 _4243_ (.A(_0567_),
    .B(_0568_),
    .ZN(_0569_));
 NAND3_X1 _4244_ (.A1(\section_2.yn2[7] ),
    .A2(\section_2.yn2[6] ),
    .A3(_0569_),
    .ZN(_0570_));
 INV_X1 _4245_ (.A(_0565_),
    .ZN(_0571_));
 NAND2_X1 _4246_ (.A1(_0563_),
    .A2(_0562_),
    .ZN(_0572_));
 XOR2_X1 _4247_ (.A(_0572_),
    .B(_0557_),
    .Z(_0573_));
 NOR2_X1 _4248_ (.A1(_0571_),
    .A2(_0573_),
    .ZN(_0574_));
 OAI21_X1 _4249_ (.A(_0568_),
    .B1(_0574_),
    .B2(_0564_),
    .ZN(_0575_));
 AOI21_X1 _4250_ (.A(_0556_),
    .B1(_0570_),
    .B2(_0575_),
    .ZN(_0576_));
 INV_X1 _4251_ (.A(\section_2.yn2[1] ),
    .ZN(_0577_));
 INV_X1 _4252_ (.A(\section_2.yn2[0] ),
    .ZN(_0578_));
 NAND2_X1 _4253_ (.A1(\section_2.yn2[3] ),
    .A2(_0578_),
    .ZN(_0579_));
 XNOR2_X1 _4254_ (.A(_0577_),
    .B(_0579_),
    .ZN(_0580_));
 NAND2_X1 _4255_ (.A1(_0575_),
    .A2(_0570_),
    .ZN(_0581_));
 XNOR2_X1 _4256_ (.A(_0581_),
    .B(_0556_),
    .ZN(_0582_));
 AOI21_X1 _4257_ (.A(_0576_),
    .B1(_0580_),
    .B2(_0582_),
    .ZN(_0583_));
 OR3_X1 _4258_ (.A1(_0521_),
    .A2(_0537_),
    .A3(_0538_),
    .ZN(_0584_));
 AOI21_X1 _4259_ (.A(_0541_),
    .B1(_0542_),
    .B2(_0584_),
    .ZN(_0585_));
 NOR3_X1 _4260_ (.A1(_0554_),
    .A2(_0583_),
    .A3(_0585_),
    .ZN(_0586_));
 OAI21_X1 _4261_ (.A(_0583_),
    .B1(_0585_),
    .B2(_0554_),
    .ZN(_0587_));
 NOR2_X1 _4262_ (.A1(\section_2.yn2[1] ),
    .A2(_0579_),
    .ZN(_0588_));
 AOI21_X1 _4263_ (.A(_0586_),
    .B1(_0587_),
    .B2(_0588_),
    .ZN(_0589_));
 XNOR2_X1 _4264_ (.A(_0519_),
    .B(_0545_),
    .ZN(_0590_));
 NOR2_X1 _4265_ (.A1(_0589_),
    .A2(_0590_),
    .ZN(_0591_));
 NAND2_X1 _4266_ (.A1(_0589_),
    .A2(_0590_),
    .ZN(_0592_));
 OAI21_X1 _4267_ (.A(_0551_),
    .B1(_0553_),
    .B2(_0539_),
    .ZN(_0593_));
 NAND3_X1 _4268_ (.A1(_0584_),
    .A2(_0541_),
    .A3(_0542_),
    .ZN(_0594_));
 AOI221_X1 _4269_ (.A(_0576_),
    .B1(_0580_),
    .B2(_0582_),
    .C1(_0593_),
    .C2(_0594_),
    .ZN(_0595_));
 NOR4_X1 _4270_ (.A1(\section_2.yn2[1] ),
    .A2(_0579_),
    .A3(_0586_),
    .A4(_0595_),
    .ZN(_0596_));
 XNOR2_X1 _4271_ (.A(_0565_),
    .B(_0573_),
    .ZN(_0597_));
 XNOR2_X1 _4272_ (.A(\section_2.yn2[6] ),
    .B(\section_2.yn2[5] ),
    .ZN(_0598_));
 XOR2_X1 _4273_ (.A(_2926_),
    .B(_2927_),
    .Z(_0599_));
 NAND2_X1 _4274_ (.A1(\section_2.yn2[7] ),
    .A2(_0599_),
    .ZN(_0600_));
 XNOR2_X1 _4275_ (.A(\section_2.yn2[7] ),
    .B(_0599_),
    .ZN(_0601_));
 OAI21_X1 _4276_ (.A(_0600_),
    .B1(_0601_),
    .B2(_0297_),
    .ZN(_0602_));
 INV_X1 _4277_ (.A(_0602_),
    .ZN(_0603_));
 XOR2_X1 _4278_ (.A(\section_2.yn2[7] ),
    .B(_0560_),
    .Z(_0604_));
 XNOR2_X1 _4279_ (.A(_0603_),
    .B(_0604_),
    .ZN(_0605_));
 NOR2_X1 _4280_ (.A1(_0598_),
    .A2(_0605_),
    .ZN(_0606_));
 NOR2_X1 _4281_ (.A1(_0603_),
    .A2(_0604_),
    .ZN(_0607_));
 OAI21_X1 _4282_ (.A(_0597_),
    .B1(_0606_),
    .B2(_0607_),
    .ZN(_0608_));
 NAND2_X1 _4283_ (.A1(\section_2.yn2[6] ),
    .A2(\section_2.yn2[5] ),
    .ZN(_0609_));
 XNOR2_X1 _4284_ (.A(_0025_),
    .B(_0609_),
    .ZN(_0610_));
 NOR2_X1 _4285_ (.A1(_0607_),
    .A2(_0606_),
    .ZN(_0611_));
 XOR2_X1 _4286_ (.A(_0611_),
    .B(_0597_),
    .Z(_0612_));
 OAI21_X1 _4287_ (.A(_0608_),
    .B1(_0610_),
    .B2(_0612_),
    .ZN(_0613_));
 NAND2_X1 _4288_ (.A1(\section_2.yn2[7] ),
    .A2(\section_2.yn2[6] ),
    .ZN(_0614_));
 XNOR2_X1 _4289_ (.A(_0614_),
    .B(_0569_),
    .ZN(_0615_));
 NAND2_X1 _4290_ (.A1(_0613_),
    .A2(_0615_),
    .ZN(_0616_));
 XOR2_X1 _4291_ (.A(\section_2.yn2[3] ),
    .B(\section_2.yn2[0] ),
    .Z(_0617_));
 OAI21_X1 _4292_ (.A(_0617_),
    .B1(_0609_),
    .B2(_0025_),
    .ZN(_0618_));
 OR3_X1 _4293_ (.A1(_0025_),
    .A2(_0609_),
    .A3(_0617_),
    .ZN(_0619_));
 NAND2_X1 _4294_ (.A1(_0618_),
    .A2(_0619_),
    .ZN(_0620_));
 XNOR2_X1 _4295_ (.A(_0613_),
    .B(_0615_),
    .ZN(_0621_));
 OAI21_X1 _4296_ (.A(_0616_),
    .B1(_0620_),
    .B2(_0621_),
    .ZN(_0622_));
 XOR2_X1 _4297_ (.A(_0580_),
    .B(_0582_),
    .Z(_0623_));
 AND2_X1 _4298_ (.A1(_0622_),
    .A2(_0623_),
    .ZN(_0624_));
 XOR2_X1 _4299_ (.A(_0622_),
    .B(_0623_),
    .Z(_0625_));
 INV_X1 _4300_ (.A(_0619_),
    .ZN(_0626_));
 AOI21_X1 _4301_ (.A(_0624_),
    .B1(_0625_),
    .B2(_0626_),
    .ZN(_0627_));
 OR3_X1 _4302_ (.A1(_0554_),
    .A2(_0583_),
    .A3(_0585_),
    .ZN(_0628_));
 AOI21_X1 _4303_ (.A(_0588_),
    .B1(_0628_),
    .B2(_0587_),
    .ZN(_0629_));
 NOR3_X1 _4304_ (.A1(_0596_),
    .A2(_0627_),
    .A3(_0629_),
    .ZN(_0630_));
 NAND2_X1 _4305_ (.A1(\section_2.yn2[5] ),
    .A2(\section_2.yn2[4] ),
    .ZN(_0631_));
 XOR2_X1 _4306_ (.A(_0027_),
    .B(_0631_),
    .Z(_0632_));
 XNOR2_X1 _4307_ (.A(_2924_),
    .B(_2925_),
    .ZN(_0633_));
 XNOR2_X1 _4308_ (.A(_0297_),
    .B(_0633_),
    .ZN(_0634_));
 OAI22_X1 _4309_ (.A1(_0026_),
    .A2(_0633_),
    .B1(_0634_),
    .B2(_0429_),
    .ZN(_0635_));
 XNOR2_X1 _4310_ (.A(_0297_),
    .B(_0601_),
    .ZN(_0636_));
 INV_X1 _4311_ (.A(_0636_),
    .ZN(_0637_));
 NAND2_X1 _4312_ (.A1(_0635_),
    .A2(_0637_),
    .ZN(_0638_));
 XNOR2_X1 _4313_ (.A(\section_2.yn2[5] ),
    .B(\section_2.yn2[4] ),
    .ZN(_0639_));
 XOR2_X1 _4314_ (.A(_0635_),
    .B(_0636_),
    .Z(_0640_));
 OAI21_X1 _4315_ (.A(_0638_),
    .B1(_0639_),
    .B2(_0640_),
    .ZN(_0641_));
 XOR2_X1 _4316_ (.A(_0598_),
    .B(_0605_),
    .Z(_0642_));
 XOR2_X1 _4317_ (.A(_0641_),
    .B(_0642_),
    .Z(_0643_));
 AND2_X1 _4318_ (.A1(_0632_),
    .A2(_0643_),
    .ZN(_0644_));
 AOI21_X1 _4319_ (.A(_0644_),
    .B1(_0642_),
    .B2(_0641_),
    .ZN(_0645_));
 XNOR2_X1 _4320_ (.A(_0610_),
    .B(_0612_),
    .ZN(_0646_));
 OR2_X1 _4321_ (.A1(_0645_),
    .A2(_0646_),
    .ZN(_0647_));
 INV_X1 _4322_ (.A(_0647_),
    .ZN(_0648_));
 XNOR2_X1 _4323_ (.A(_0645_),
    .B(_0646_),
    .ZN(_0649_));
 NOR3_X1 _4324_ (.A1(_0027_),
    .A2(_0631_),
    .A3(_0649_),
    .ZN(_0650_));
 NOR2_X1 _4325_ (.A1(_0648_),
    .A2(_0650_),
    .ZN(_0651_));
 XNOR2_X1 _4326_ (.A(_0620_),
    .B(_0621_),
    .ZN(_0652_));
 OR2_X1 _4327_ (.A1(_0651_),
    .A2(_0652_),
    .ZN(_0653_));
 INV_X1 _4328_ (.A(_0653_),
    .ZN(_0654_));
 XNOR2_X1 _4329_ (.A(_0619_),
    .B(_0625_),
    .ZN(_0655_));
 NAND2_X1 _4330_ (.A1(_0654_),
    .A2(_0655_),
    .ZN(_0656_));
 XNOR2_X1 _4331_ (.A(_0654_),
    .B(_0655_),
    .ZN(_0657_));
 NOR2_X1 _4332_ (.A1(_0027_),
    .A2(_0631_),
    .ZN(_0658_));
 XNOR2_X1 _4333_ (.A(_0658_),
    .B(_0649_),
    .ZN(_0659_));
 NAND2_X1 _4334_ (.A1(\section_2.yn2[4] ),
    .A2(\section_2.yn2[3] ),
    .ZN(_0660_));
 NOR2_X1 _4335_ (.A1(_0029_),
    .A2(_0660_),
    .ZN(_0661_));
 XNOR2_X1 _4336_ (.A(_0632_),
    .B(_0643_),
    .ZN(_0662_));
 XOR2_X1 _4337_ (.A(_0029_),
    .B(_0660_),
    .Z(_0663_));
 XNOR2_X1 _4338_ (.A(_2922_),
    .B(_2923_),
    .ZN(_0664_));
 XNOR2_X1 _4339_ (.A(_0429_),
    .B(_0664_),
    .ZN(_0665_));
 OAI22_X1 _4340_ (.A1(_0028_),
    .A2(_0664_),
    .B1(_0665_),
    .B2(_0516_),
    .ZN(_0666_));
 XNOR2_X1 _4341_ (.A(\section_2.yn2[5] ),
    .B(_0634_),
    .ZN(_0667_));
 NAND2_X1 _4342_ (.A1(_0666_),
    .A2(_0667_),
    .ZN(_0668_));
 XNOR2_X1 _4343_ (.A(\section_2.yn2[4] ),
    .B(\section_2.yn2[3] ),
    .ZN(_0669_));
 XNOR2_X1 _4344_ (.A(_0666_),
    .B(_0667_),
    .ZN(_0670_));
 OAI21_X1 _4345_ (.A(_0668_),
    .B1(_0669_),
    .B2(_0670_),
    .ZN(_0671_));
 XOR2_X1 _4346_ (.A(_0639_),
    .B(_0640_),
    .Z(_0672_));
 XNOR2_X1 _4347_ (.A(_0671_),
    .B(_0672_),
    .ZN(_0673_));
 INV_X1 _4348_ (.A(_0673_),
    .ZN(_0674_));
 NAND2_X1 _4349_ (.A1(_0663_),
    .A2(_0674_),
    .ZN(_0675_));
 NAND2_X1 _4350_ (.A1(_0671_),
    .A2(_0672_),
    .ZN(_0676_));
 AOI21_X1 _4351_ (.A(_0662_),
    .B1(_0675_),
    .B2(_0676_),
    .ZN(_0677_));
 AND3_X1 _4352_ (.A1(_0676_),
    .A2(_0675_),
    .A3(_0662_),
    .ZN(_0678_));
 NOR2_X1 _4353_ (.A1(_0677_),
    .A2(_0678_),
    .ZN(_0679_));
 AND2_X1 _4354_ (.A1(_0661_),
    .A2(_0679_),
    .ZN(_0680_));
 OAI21_X1 _4355_ (.A(_0659_),
    .B1(_0680_),
    .B2(_0677_),
    .ZN(_0681_));
 XNOR2_X1 _4356_ (.A(_0651_),
    .B(_0652_),
    .ZN(_0682_));
 NOR2_X1 _4357_ (.A1(_0681_),
    .A2(_0682_),
    .ZN(_0683_));
 OR3_X1 _4358_ (.A1(_0677_),
    .A2(_0680_),
    .A3(_0659_),
    .ZN(_0684_));
 NAND2_X1 _4359_ (.A1(_0681_),
    .A2(_0684_),
    .ZN(_0685_));
 NOR2_X1 _4360_ (.A1(_0661_),
    .A2(_0679_),
    .ZN(_0686_));
 XOR2_X1 _4361_ (.A(_0669_),
    .B(_0670_),
    .Z(_0687_));
 XNOR2_X1 _4362_ (.A(\section_2.yn2[3] ),
    .B(\section_2.yn2[2] ),
    .ZN(_0688_));
 XOR2_X1 _4363_ (.A(_2920_),
    .B(_2921_),
    .Z(_0689_));
 NAND2_X1 _4364_ (.A1(\section_2.yn2[4] ),
    .A2(_0689_),
    .ZN(_0690_));
 XNOR2_X1 _4365_ (.A(\section_2.yn2[4] ),
    .B(_0689_),
    .ZN(_0691_));
 OAI21_X1 _4366_ (.A(_0690_),
    .B1(_0691_),
    .B2(_0498_),
    .ZN(_0692_));
 XNOR2_X1 _4367_ (.A(\section_2.yn2[4] ),
    .B(_0665_),
    .ZN(_0693_));
 XNOR2_X1 _4368_ (.A(_0692_),
    .B(_0693_),
    .ZN(_0694_));
 NOR2_X1 _4369_ (.A1(_0688_),
    .A2(_0694_),
    .ZN(_0695_));
 AND2_X1 _4370_ (.A1(_0692_),
    .A2(_0693_),
    .ZN(_0696_));
 OAI21_X1 _4371_ (.A(_0687_),
    .B1(_0695_),
    .B2(_0696_),
    .ZN(_0697_));
 OR3_X1 _4372_ (.A1(_0696_),
    .A2(_0695_),
    .A3(_0687_),
    .ZN(_0698_));
 NAND2_X1 _4373_ (.A1(_0697_),
    .A2(_0698_),
    .ZN(_0699_));
 NAND2_X1 _4374_ (.A1(\section_2.yn2[3] ),
    .A2(\section_2.yn2[2] ),
    .ZN(_0700_));
 OAI21_X1 _4375_ (.A(_0697_),
    .B1(_0699_),
    .B2(_0700_),
    .ZN(_0701_));
 XNOR2_X1 _4376_ (.A(_0663_),
    .B(_0673_),
    .ZN(_0702_));
 NAND2_X1 _4377_ (.A1(_0701_),
    .A2(_0702_),
    .ZN(_0703_));
 OR3_X1 _4378_ (.A1(_0680_),
    .A2(_0686_),
    .A3(_0703_),
    .ZN(_0704_));
 OAI21_X1 _4379_ (.A(_0703_),
    .B1(_0686_),
    .B2(_0680_),
    .ZN(_0705_));
 NOR2_X1 _4380_ (.A1(_0700_),
    .A2(_0699_),
    .ZN(_0706_));
 XNOR2_X1 _4381_ (.A(_0688_),
    .B(_0694_),
    .ZN(_0707_));
 XOR2_X1 _4382_ (.A(\section_2.yn2[2] ),
    .B(\section_2.yn2[1] ),
    .Z(_0708_));
 XNOR2_X1 _4383_ (.A(_2862_),
    .B(_2919_),
    .ZN(_0709_));
 NOR2_X1 _4384_ (.A1(_0498_),
    .A2(_0709_),
    .ZN(_0710_));
 XNOR2_X1 _4385_ (.A(_0498_),
    .B(_0709_),
    .ZN(_0711_));
 NOR2_X1 _4386_ (.A1(_0540_),
    .A2(_0711_),
    .ZN(_0712_));
 NOR2_X1 _4387_ (.A1(_0710_),
    .A2(_0712_),
    .ZN(_0713_));
 XNOR2_X1 _4388_ (.A(_0498_),
    .B(_0691_),
    .ZN(_0714_));
 XOR2_X1 _4389_ (.A(_0713_),
    .B(_0714_),
    .Z(_0715_));
 NAND2_X1 _4390_ (.A1(_0708_),
    .A2(_0715_),
    .ZN(_0716_));
 OR2_X1 _4391_ (.A1(_0713_),
    .A2(_0714_),
    .ZN(_0717_));
 AOI21_X1 _4392_ (.A(_0707_),
    .B1(_0716_),
    .B2(_0717_),
    .ZN(_0718_));
 AND3_X1 _4393_ (.A1(_0717_),
    .A2(_0716_),
    .A3(_0707_),
    .ZN(_0719_));
 NOR2_X1 _4394_ (.A1(_0718_),
    .A2(_0719_),
    .ZN(_0720_));
 AND3_X1 _4395_ (.A1(\section_2.yn2[2] ),
    .A2(\section_2.yn2[1] ),
    .A3(_0720_),
    .ZN(_0721_));
 NOR2_X1 _4396_ (.A1(_0718_),
    .A2(_0721_),
    .ZN(_0722_));
 AND2_X1 _4397_ (.A1(_0700_),
    .A2(_0699_),
    .ZN(_0723_));
 OR3_X1 _4398_ (.A1(_0706_),
    .A2(_0722_),
    .A3(_0723_),
    .ZN(_0724_));
 XNOR2_X1 _4399_ (.A(_0701_),
    .B(_0702_),
    .ZN(_0725_));
 NAND2_X1 _4400_ (.A1(_0724_),
    .A2(_0725_),
    .ZN(_0726_));
 OAI21_X1 _4401_ (.A(_0722_),
    .B1(_0723_),
    .B2(_0706_),
    .ZN(_0727_));
 NAND2_X1 _4402_ (.A1(_0724_),
    .A2(_0727_),
    .ZN(_0728_));
 XNOR2_X1 _4403_ (.A(_0708_),
    .B(_0715_),
    .ZN(_0729_));
 NOR2_X1 _4404_ (.A1(\section_2.yn2[1] ),
    .A2(\section_2.yn2[0] ),
    .ZN(_0730_));
 NOR2_X1 _4405_ (.A1(_0577_),
    .A2(_0578_),
    .ZN(_0731_));
 NAND2_X1 _4406_ (.A1(\section_2.xn2[0] ),
    .A2(_2409_),
    .ZN(_0732_));
 XOR2_X1 _4407_ (.A(_2394_),
    .B(_0732_),
    .Z(_0733_));
 XNOR2_X1 _4408_ (.A(_0540_),
    .B(_0733_),
    .ZN(_0734_));
 OAI22_X1 _4409_ (.A1(_0025_),
    .A2(_0733_),
    .B1(_0734_),
    .B2(_0577_),
    .ZN(_0735_));
 XNOR2_X1 _4410_ (.A(_0540_),
    .B(_0711_),
    .ZN(_0736_));
 XOR2_X1 _4411_ (.A(_0735_),
    .B(_0736_),
    .Z(_0737_));
 OR3_X1 _4412_ (.A1(_0730_),
    .A2(_0731_),
    .A3(_0737_),
    .ZN(_0738_));
 INV_X1 _4413_ (.A(_0736_),
    .ZN(_0739_));
 NAND2_X1 _4414_ (.A1(_0735_),
    .A2(_0739_),
    .ZN(_0740_));
 AOI21_X1 _4415_ (.A(_0729_),
    .B1(_0738_),
    .B2(_0740_),
    .ZN(_0741_));
 NAND2_X1 _4416_ (.A1(_0740_),
    .A2(_0738_),
    .ZN(_0742_));
 XNOR2_X1 _4417_ (.A(_0742_),
    .B(_0729_),
    .ZN(_0743_));
 AOI21_X1 _4418_ (.A(_0741_),
    .B1(_0743_),
    .B2(_0731_),
    .ZN(_0744_));
 AOI21_X1 _4419_ (.A(_0720_),
    .B1(\section_2.yn2[1] ),
    .B2(\section_2.yn2[2] ),
    .ZN(_0745_));
 NOR3_X1 _4420_ (.A1(_0721_),
    .A2(_0744_),
    .A3(_0745_),
    .ZN(_0746_));
 OAI21_X1 _4421_ (.A(_0744_),
    .B1(_0745_),
    .B2(_0721_),
    .ZN(_0747_));
 XNOR2_X1 _4422_ (.A(_0731_),
    .B(_0743_),
    .ZN(_0748_));
 INV_X1 _4423_ (.A(\coll_reg[0] ),
    .ZN(_0749_));
 NAND2_X1 _4424_ (.A1(_0749_),
    .A2(\section_2.xn2[0] ),
    .ZN(_0750_));
 NAND2_X1 _4425_ (.A1(\coll_reg[0] ),
    .A2(_2390_),
    .ZN(_0751_));
 AOI21_X1 _4426_ (.A(_0029_),
    .B1(_0750_),
    .B2(_0751_),
    .ZN(_0752_));
 XNOR2_X1 _4427_ (.A(_2389_),
    .B(_0750_),
    .ZN(_0753_));
 XNOR2_X1 _4428_ (.A(_0577_),
    .B(_0753_),
    .ZN(_0754_));
 OAI22_X1 _4429_ (.A1(_0027_),
    .A2(_0753_),
    .B1(_0754_),
    .B2(_0578_),
    .ZN(_0755_));
 XNOR2_X1 _4430_ (.A(_0577_),
    .B(_0734_),
    .ZN(_0756_));
 XNOR2_X1 _4431_ (.A(_0755_),
    .B(_0756_),
    .ZN(_0757_));
 NAND2_X1 _4432_ (.A1(\section_2.yn2[0] ),
    .A2(_0757_),
    .ZN(_0758_));
 OAI21_X1 _4433_ (.A(_0737_),
    .B1(_0731_),
    .B2(_0730_),
    .ZN(_0759_));
 INV_X1 _4434_ (.A(_0755_),
    .ZN(_0760_));
 OAI21_X1 _4435_ (.A(_0758_),
    .B1(_0756_),
    .B2(_0760_),
    .ZN(_0761_));
 NAND3_X1 _4436_ (.A1(_0738_),
    .A2(_0759_),
    .A3(_0761_),
    .ZN(_0762_));
 NOR2_X1 _4437_ (.A1(_0754_),
    .A2(_0757_),
    .ZN(_0763_));
 AOI21_X1 _4438_ (.A(_0761_),
    .B1(_0759_),
    .B2(_0738_),
    .ZN(_0764_));
 AOI211_X1 _4439_ (.A(_0763_),
    .B(_0764_),
    .C1(_0578_),
    .C2(_0754_),
    .ZN(_0765_));
 NAND4_X1 _4440_ (.A1(_0752_),
    .A2(_0758_),
    .A3(_0762_),
    .A4(_0765_),
    .ZN(_0766_));
 AOI21_X1 _4441_ (.A(_0748_),
    .B1(_0766_),
    .B2(_0762_),
    .ZN(_0767_));
 AOI21_X1 _4442_ (.A(_0746_),
    .B1(_0747_),
    .B2(_0767_),
    .ZN(_0768_));
 OAI22_X1 _4443_ (.A1(_0724_),
    .A2(_0725_),
    .B1(_0728_),
    .B2(_0768_),
    .ZN(_0769_));
 NAND3_X1 _4444_ (.A1(_0705_),
    .A2(_0726_),
    .A3(_0769_),
    .ZN(_0770_));
 AOI21_X1 _4445_ (.A(_0685_),
    .B1(_0704_),
    .B2(_0770_),
    .ZN(_0771_));
 XOR2_X1 _4446_ (.A(_0681_),
    .B(_0682_),
    .Z(_0772_));
 AOI21_X1 _4447_ (.A(_0683_),
    .B1(_0771_),
    .B2(_0772_),
    .ZN(_0773_));
 OAI21_X1 _4448_ (.A(_0656_),
    .B1(_0657_),
    .B2(_0773_),
    .ZN(_0774_));
 XNOR2_X1 _4449_ (.A(_0589_),
    .B(_0590_),
    .ZN(_0775_));
 OAI22_X1 _4450_ (.A1(\section_2.yn2[1] ),
    .A2(_0579_),
    .B1(_0586_),
    .B2(_0595_),
    .ZN(_0776_));
 NAND3_X1 _4451_ (.A1(_0588_),
    .A2(_0628_),
    .A3(_0587_),
    .ZN(_0777_));
 AOI221_X1 _4452_ (.A(_0624_),
    .B1(_0625_),
    .B2(_0626_),
    .C1(_0776_),
    .C2(_0777_),
    .ZN(_0778_));
 NOR3_X1 _4453_ (.A1(_0775_),
    .A2(_0630_),
    .A3(_0778_),
    .ZN(_0779_));
 AOI221_X1 _4454_ (.A(_0591_),
    .B1(_0592_),
    .B2(_0630_),
    .C1(_0774_),
    .C2(_0779_),
    .ZN(_0780_));
 OAI21_X1 _4455_ (.A(_0548_),
    .B1(_0550_),
    .B2(_0780_),
    .ZN(_0781_));
 AOI21_X1 _4456_ (.A(_0513_),
    .B1(_0514_),
    .B2(_0781_),
    .ZN(_0782_));
 OAI21_X1 _4457_ (.A(_0475_),
    .B1(_0477_),
    .B2(_0782_),
    .ZN(_0783_));
 XOR2_X1 _4458_ (.A(_0365_),
    .B(_0418_),
    .Z(_0784_));
 AOI21_X1 _4459_ (.A(_0419_),
    .B1(_0783_),
    .B2(_0784_),
    .ZN(_0785_));
 OR2_X1 _4460_ (.A1(_0368_),
    .A2(_0416_),
    .ZN(_0786_));
 OAI21_X1 _4461_ (.A(_0786_),
    .B1(_0417_),
    .B2(_0366_),
    .ZN(_0787_));
 NOR2_X1 _4462_ (.A1(_0442_),
    .A2(\section_2.yn2[8] ),
    .ZN(_0788_));
 NOR3_X1 _4463_ (.A1(_0293_),
    .A2(_0369_),
    .A3(_0413_),
    .ZN(_0789_));
 OR2_X1 _4464_ (.A1(_0370_),
    .A2(_0414_),
    .ZN(_0790_));
 INV_X1 _4465_ (.A(_1264_),
    .ZN(_0791_));
 AOI21_X1 _4466_ (.A(_0789_),
    .B1(_0790_),
    .B2(_0791_),
    .ZN(_0792_));
 NOR3_X1 _4467_ (.A1(_0002_),
    .A2(_0358_),
    .A3(_0413_),
    .ZN(_0793_));
 OAI21_X1 _4468_ (.A(_0442_),
    .B1(_0410_),
    .B2(_0411_),
    .ZN(_0794_));
 OR3_X1 _4469_ (.A1(_0442_),
    .A2(_0410_),
    .A3(_0411_),
    .ZN(_0795_));
 AOI21_X1 _4470_ (.A(_0002_),
    .B1(_0794_),
    .B2(_0795_),
    .ZN(_0796_));
 NOR2_X1 _4471_ (.A1(_0348_),
    .A2(_0407_),
    .ZN(_0797_));
 AOI21_X1 _4472_ (.A(_0797_),
    .B1(_0408_),
    .B2(_0371_),
    .ZN(_0798_));
 NAND2_X1 _4473_ (.A1(_0350_),
    .A2(_0408_),
    .ZN(_0799_));
 NAND4_X1 _4474_ (.A1(_0219_),
    .A2(_0291_),
    .A3(_0350_),
    .A4(_0408_),
    .ZN(_0800_));
 NOR2_X1 _4475_ (.A1(_2861_),
    .A2(_0168_),
    .ZN(_0801_));
 OAI21_X1 _4476_ (.A(_0448_),
    .B1(_2894_),
    .B2(_0446_),
    .ZN(_0802_));
 AOI221_X1 _4477_ (.A(_0220_),
    .B1(_0221_),
    .B2(_0222_),
    .C1(_0801_),
    .C2(_0802_),
    .ZN(_0803_));
 OAI221_X1 _4478_ (.A(_0798_),
    .B1(_0799_),
    .B2(_0354_),
    .C1(_0800_),
    .C2(_0803_),
    .ZN(_0804_));
 NOR3_X1 _4479_ (.A1(_0446_),
    .A2(_2881_),
    .A3(_2932_),
    .ZN(_0805_));
 NAND2_X1 _4480_ (.A1(_0805_),
    .A2(_0801_),
    .ZN(_0806_));
 NOR3_X1 _4481_ (.A1(_2931_),
    .A2(_0806_),
    .A3(_0800_),
    .ZN(_0807_));
 NOR2_X1 _4482_ (.A1(_0804_),
    .A2(_0807_),
    .ZN(_0808_));
 AND2_X1 _4483_ (.A1(_0377_),
    .A2(_0406_),
    .ZN(_0809_));
 NOR2_X1 _4484_ (.A1(z[9]),
    .A2(_0316_),
    .ZN(_0810_));
 NAND2_X1 _4485_ (.A1(_0382_),
    .A2(_0403_),
    .ZN(_0811_));
 NAND2_X1 _4486_ (.A1(z[10]),
    .A2(_0402_),
    .ZN(_0812_));
 INV_X1 _4487_ (.A(_0812_),
    .ZN(_0813_));
 NAND2_X1 _4488_ (.A1(_0342_),
    .A2(_0813_),
    .ZN(_0814_));
 OAI21_X1 _4489_ (.A(_0811_),
    .B1(_0814_),
    .B2(_0285_),
    .ZN(_0815_));
 NOR2_X1 _4490_ (.A1(_2767_),
    .A2(z[8]),
    .ZN(_0816_));
 XNOR2_X1 _4491_ (.A(_2951_),
    .B(_0816_),
    .ZN(_0817_));
 OR2_X1 _4492_ (.A1(_0386_),
    .A2(_0400_),
    .ZN(_0818_));
 OAI21_X1 _4493_ (.A(_0818_),
    .B1(_0401_),
    .B2(_0384_),
    .ZN(_0819_));
 MUX2_X1 _4494_ (.A(_0396_),
    .B(_0031_),
    .S(_0394_),
    .Z(_0820_));
 MUX2_X1 _4495_ (.A(_0395_),
    .B(_0398_),
    .S(\section_2.xn2[10] ),
    .Z(_0821_));
 XNOR2_X1 _4496_ (.A(_0820_),
    .B(_0821_),
    .ZN(_0822_));
 XNOR2_X1 _4497_ (.A(_0819_),
    .B(_0822_),
    .ZN(_0823_));
 AOI21_X1 _4498_ (.A(_0823_),
    .B1(_0813_),
    .B2(_0342_),
    .ZN(_0824_));
 XNOR2_X1 _4499_ (.A(_0817_),
    .B(_0824_),
    .ZN(_0825_));
 XNOR2_X1 _4500_ (.A(_0815_),
    .B(_0825_),
    .ZN(_0826_));
 XNOR2_X1 _4501_ (.A(_0810_),
    .B(_0826_),
    .ZN(_0827_));
 NOR3_X1 _4502_ (.A1(z[8]),
    .A2(_0243_),
    .A3(_0405_),
    .ZN(_0828_));
 INV_X1 _4503_ (.A(_0404_),
    .ZN(_0829_));
 NOR2_X1 _4504_ (.A1(_0380_),
    .A2(_0829_),
    .ZN(_0830_));
 OAI21_X1 _4505_ (.A(_0827_),
    .B1(_0828_),
    .B2(_0830_),
    .ZN(_0831_));
 OR3_X1 _4506_ (.A1(_0830_),
    .A2(_0828_),
    .A3(_0827_),
    .ZN(_0832_));
 NAND2_X1 _4507_ (.A1(_0831_),
    .A2(_0832_),
    .ZN(_0833_));
 XNOR2_X1 _4508_ (.A(_0809_),
    .B(_0833_),
    .ZN(_0834_));
 XNOR2_X1 _4509_ (.A(_0808_),
    .B(_0834_),
    .ZN(_0835_));
 XNOR2_X1 _4510_ (.A(\section_2.yn2[10] ),
    .B(_0835_),
    .ZN(_0836_));
 XNOR2_X1 _4511_ (.A(_0796_),
    .B(_0836_),
    .ZN(_0837_));
 XNOR2_X1 _4512_ (.A(_0793_),
    .B(_0837_),
    .ZN(_0838_));
 XNOR2_X1 _4513_ (.A(_0458_),
    .B(_0838_),
    .ZN(_0839_));
 XNOR2_X1 _4514_ (.A(_0792_),
    .B(_0839_),
    .ZN(_0840_));
 XOR2_X1 _4515_ (.A(_0788_),
    .B(_0840_),
    .Z(_0841_));
 XOR2_X1 _4516_ (.A(_0787_),
    .B(_0841_),
    .Z(_0842_));
 XOR2_X1 _4517_ (.A(_0785_),
    .B(_0842_),
    .Z(_0843_));
 XNOR2_X1 _4518_ (.A(_0783_),
    .B(_0784_),
    .ZN(_0844_));
 OR2_X1 _4519_ (.A1(_0472_),
    .A2(_0473_),
    .ZN(_0845_));
 INV_X1 _4520_ (.A(_0476_),
    .ZN(_0846_));
 OAI21_X1 _4521_ (.A(_0845_),
    .B1(_0782_),
    .B2(_0846_),
    .ZN(_0847_));
 XNOR2_X1 _4522_ (.A(_0441_),
    .B(_0847_),
    .ZN(_0848_));
 XNOR2_X1 _4523_ (.A(_0782_),
    .B(_0476_),
    .ZN(_0849_));
 XOR2_X1 _4524_ (.A(_0514_),
    .B(_0781_),
    .Z(_0850_));
 XNOR2_X1 _4525_ (.A(_0550_),
    .B(_0780_),
    .ZN(_0851_));
 NOR2_X1 _4526_ (.A1(_0630_),
    .A2(_0778_),
    .ZN(_0852_));
 XOR2_X1 _4527_ (.A(_0852_),
    .B(_0774_),
    .Z(_0853_));
 NAND3_X1 _4528_ (.A1(_0685_),
    .A2(_0704_),
    .A3(_0770_),
    .ZN(_0854_));
 NAND2_X1 _4529_ (.A1(_0772_),
    .A2(_0854_),
    .ZN(_0855_));
 NOR2_X1 _4530_ (.A1(_0771_),
    .A2(_0855_),
    .ZN(_0856_));
 XOR2_X1 _4531_ (.A(_0657_),
    .B(_0773_),
    .Z(_0857_));
 AND2_X1 _4532_ (.A1(_0856_),
    .A2(_0857_),
    .ZN(_0858_));
 AND2_X1 _4533_ (.A1(_0853_),
    .A2(_0858_),
    .ZN(_0859_));
 AOI21_X1 _4534_ (.A(_0630_),
    .B1(_0852_),
    .B2(_0774_),
    .ZN(_0860_));
 XOR2_X1 _4535_ (.A(_0775_),
    .B(_0860_),
    .Z(_0861_));
 NAND2_X1 _4536_ (.A1(_0859_),
    .A2(_0861_),
    .ZN(_0862_));
 NOR2_X1 _4537_ (.A1(_0851_),
    .A2(_0862_),
    .ZN(_0863_));
 NAND3_X1 _4538_ (.A1(_0849_),
    .A2(_0850_),
    .A3(_0863_),
    .ZN(_0864_));
 OR3_X1 _4539_ (.A1(_0844_),
    .A2(_0848_),
    .A3(_0864_),
    .ZN(_0865_));
 OAI21_X1 _4540_ (.A(_1253_),
    .B1(_0843_),
    .B2(_0865_),
    .ZN(_0866_));
 AOI21_X1 _4541_ (.A(_0866_),
    .B1(_0865_),
    .B2(_0843_),
    .ZN(_0119_));
 NAND2_X1 _4542_ (.A1(_1253_),
    .A2(_0865_),
    .ZN(_0867_));
 OR2_X1 _4543_ (.A1(_0848_),
    .A2(_0864_),
    .ZN(_0868_));
 AOI21_X1 _4544_ (.A(_0867_),
    .B1(_0868_),
    .B2(_0844_),
    .ZN(_0118_));
 NAND2_X1 _4545_ (.A1(_1253_),
    .A2(_0868_),
    .ZN(_0869_));
 AOI21_X1 _4546_ (.A(_0869_),
    .B1(_0864_),
    .B2(_0848_),
    .ZN(_0117_));
 AOI21_X1 _4547_ (.A(_0849_),
    .B1(_0850_),
    .B2(_0863_),
    .ZN(_0870_));
 NAND2_X1 _4548_ (.A1(_1253_),
    .A2(_0864_),
    .ZN(_0871_));
 NOR2_X1 _4549_ (.A1(_0870_),
    .A2(_0871_),
    .ZN(_0116_));
 OAI21_X1 _4550_ (.A(_1253_),
    .B1(_0850_),
    .B2(_0863_),
    .ZN(_0872_));
 AOI21_X1 _4551_ (.A(_0872_),
    .B1(_0863_),
    .B2(_0850_),
    .ZN(_0115_));
 AND2_X1 _4552_ (.A1(_0851_),
    .A2(_0862_),
    .ZN(_0873_));
 NOR3_X1 _4553_ (.A1(rst),
    .A2(_0863_),
    .A3(_0873_),
    .ZN(_0114_));
 OAI21_X1 _4554_ (.A(_1253_),
    .B1(_0859_),
    .B2(_0861_),
    .ZN(_0874_));
 AOI21_X1 _4555_ (.A(_0874_),
    .B1(_0861_),
    .B2(_0859_),
    .ZN(_0113_));
 NOR2_X1 _4556_ (.A1(_0853_),
    .A2(_0858_),
    .ZN(_0875_));
 NOR3_X1 _4557_ (.A1(rst),
    .A2(_0859_),
    .A3(_0875_),
    .ZN(_0112_));
 NOR2_X1 _4558_ (.A1(_0856_),
    .A2(_0857_),
    .ZN(_0876_));
 NOR3_X1 _4559_ (.A1(rst),
    .A2(_0858_),
    .A3(_0876_),
    .ZN(_0111_));
 NAND2_X1 _4560_ (.A1(_0787_),
    .A2(_0841_),
    .ZN(_0877_));
 NAND2_X1 _4561_ (.A1(_0419_),
    .A2(_0842_),
    .ZN(_0878_));
 NAND2_X1 _4562_ (.A1(_0784_),
    .A2(_0842_),
    .ZN(_0879_));
 OAI211_X1 _4563_ (.A(_0877_),
    .B(_0878_),
    .C1(_0879_),
    .C2(_0475_),
    .ZN(_0880_));
 NOR3_X1 _4564_ (.A1(_0782_),
    .A2(_0477_),
    .A3(_0879_),
    .ZN(_0881_));
 NOR2_X1 _4565_ (.A1(_0880_),
    .A2(_0881_),
    .ZN(_0882_));
 NOR2_X1 _4566_ (.A1(_1264_),
    .A2(_0415_),
    .ZN(_0883_));
 OAI21_X1 _4567_ (.A(_0839_),
    .B1(_0883_),
    .B2(_0789_),
    .ZN(_0884_));
 INV_X1 _4568_ (.A(_0884_),
    .ZN(_0885_));
 AOI21_X1 _4569_ (.A(_0885_),
    .B1(_0840_),
    .B2(_0788_),
    .ZN(_0886_));
 NOR2_X1 _4570_ (.A1(_0442_),
    .A2(\section_2.yn2[9] ),
    .ZN(_0887_));
 NAND2_X1 _4571_ (.A1(_0793_),
    .A2(_0837_),
    .ZN(_0888_));
 OAI21_X1 _4572_ (.A(_0888_),
    .B1(_0838_),
    .B2(_0231_),
    .ZN(_0889_));
 AOI211_X1 _4573_ (.A(_0002_),
    .B(_0836_),
    .C1(_0795_),
    .C2(_0794_),
    .ZN(_0890_));
 NAND3_X1 _4574_ (.A1(_0809_),
    .A2(_0831_),
    .A3(_0832_),
    .ZN(_0891_));
 INV_X1 _4575_ (.A(_0834_),
    .ZN(_0892_));
 OAI21_X1 _4576_ (.A(_0891_),
    .B1(_0892_),
    .B2(_0808_),
    .ZN(_0893_));
 NOR3_X1 _4577_ (.A1(z[9]),
    .A2(_0316_),
    .A3(_0826_),
    .ZN(_0894_));
 AOI21_X1 _4578_ (.A(_0894_),
    .B1(_0825_),
    .B2(_0815_),
    .ZN(_0895_));
 NOR3_X1 _4579_ (.A1(_0342_),
    .A2(_0812_),
    .A3(_0823_),
    .ZN(_0896_));
 OR2_X1 _4580_ (.A1(_0813_),
    .A2(_0823_),
    .ZN(_0897_));
 AOI21_X1 _4581_ (.A(_0896_),
    .B1(_0897_),
    .B2(_0817_),
    .ZN(_0898_));
 AOI21_X1 _4582_ (.A(_2767_),
    .B1(_2626_),
    .B2(_2951_),
    .ZN(_0899_));
 XNOR2_X1 _4583_ (.A(_0897_),
    .B(_0899_),
    .ZN(_0900_));
 XNOR2_X1 _4584_ (.A(_0898_),
    .B(_0900_),
    .ZN(_0901_));
 XNOR2_X1 _4585_ (.A(_0895_),
    .B(_0901_),
    .ZN(_0902_));
 XNOR2_X1 _4586_ (.A(_0831_),
    .B(_0902_),
    .ZN(_0903_));
 XNOR2_X1 _4587_ (.A(_0893_),
    .B(_0903_),
    .ZN(_0904_));
 NOR2_X1 _4588_ (.A1(_0304_),
    .A2(\section_2.yn2[10] ),
    .ZN(_0905_));
 AOI21_X1 _4589_ (.A(_0905_),
    .B1(_0835_),
    .B2(_0304_),
    .ZN(_0906_));
 XNOR2_X1 _4590_ (.A(_0904_),
    .B(_0906_),
    .ZN(_0907_));
 XNOR2_X1 _4591_ (.A(_0890_),
    .B(_0907_),
    .ZN(_0908_));
 XNOR2_X1 _4592_ (.A(_0889_),
    .B(_0908_),
    .ZN(_0909_));
 XNOR2_X1 _4593_ (.A(_0887_),
    .B(_0909_),
    .ZN(_0910_));
 XNOR2_X1 _4594_ (.A(_0886_),
    .B(_0910_),
    .ZN(_0911_));
 XNOR2_X1 _4595_ (.A(_0882_),
    .B(_0911_),
    .ZN(_0912_));
 OAI21_X1 _4596_ (.A(_0912_),
    .B1(_0865_),
    .B2(_0843_),
    .ZN(_0913_));
 OR3_X1 _4597_ (.A1(_0843_),
    .A2(_0865_),
    .A3(_0912_),
    .ZN(_0914_));
 AND3_X1 _4598_ (.A1(_1253_),
    .A2(_0913_),
    .A3(_0914_),
    .ZN(_0110_));
 OR2_X1 _4599_ (.A1(_0772_),
    .A2(_0854_),
    .ZN(_0915_));
 AND3_X1 _4600_ (.A1(_1253_),
    .A2(_0855_),
    .A3(_0915_),
    .ZN(_0109_));
 NOR2_X1 _4601_ (.A1(rst),
    .A2(net70),
    .ZN(_0108_));
 NOR2_X1 _4602_ (.A1(rst),
    .A2(_2626_),
    .ZN(_0107_));
 AND2_X1 _4603_ (.A1(_1253_),
    .A2(net58),
    .ZN(_0106_));
 AND2_X1 _4604_ (.A1(_1253_),
    .A2(net75),
    .ZN(_0105_));
 AND2_X1 _4605_ (.A1(_1253_),
    .A2(net48),
    .ZN(_0104_));
 AND2_X1 _4606_ (.A1(_1253_),
    .A2(net52),
    .ZN(_0103_));
 AND2_X1 _4607_ (.A1(_1253_),
    .A2(net50),
    .ZN(_0102_));
 AND2_X1 _4608_ (.A1(_1253_),
    .A2(net56),
    .ZN(_0101_));
 AND2_X1 _4609_ (.A1(_1253_),
    .A2(net54),
    .ZN(_0100_));
 NOR2_X1 _4610_ (.A1(rst),
    .A2(_2951_),
    .ZN(_0099_));
 NOR2_X1 _4611_ (.A1(rst),
    .A2(net61),
    .ZN(_0098_));
 NOR2_X1 _4612_ (.A1(rst),
    .A2(_2572_),
    .ZN(_0097_));
 NOR2_X1 _4613_ (.A1(rst),
    .A2(net78),
    .ZN(_0096_));
 NOR2_X1 _4614_ (.A1(rst),
    .A2(_2443_),
    .ZN(_0095_));
 NOR2_X1 _4615_ (.A1(rst),
    .A2(net64),
    .ZN(_0094_));
 NOR2_X1 _4616_ (.A1(rst),
    .A2(_2275_),
    .ZN(_0093_));
 INV_X1 _4617_ (.A(net80),
    .ZN(_0916_));
 NOR2_X1 _4618_ (.A1(rst),
    .A2(_0916_),
    .ZN(_0092_));
 INV_X1 _4619_ (.A(net65),
    .ZN(_0917_));
 NOR2_X1 _4620_ (.A1(rst),
    .A2(net66),
    .ZN(_0091_));
 NOR2_X1 _4621_ (.A1(rst),
    .A2(net72),
    .ZN(_0090_));
 NOR2_X1 _4622_ (.A1(rst),
    .A2(_1330_),
    .ZN(_0089_));
 NOR2_X1 _4623_ (.A1(rst),
    .A2(_2717_),
    .ZN(_0088_));
 NOR2_X1 _4624_ (.A1(rst),
    .A2(net42),
    .ZN(_0087_));
 AND2_X1 _4625_ (.A1(_1253_),
    .A2(net67),
    .ZN(_0086_));
 NOR2_X1 _4626_ (.A1(rst),
    .A2(_2585_),
    .ZN(_0085_));
 INV_X1 _4627_ (.A(net113),
    .ZN(_0918_));
 NOR2_X1 _4628_ (.A1(rst),
    .A2(_0918_),
    .ZN(_0084_));
 AND2_X1 _4629_ (.A1(_1253_),
    .A2(net88),
    .ZN(_0083_));
 NOR2_X1 _4630_ (.A1(rst),
    .A2(_2283_),
    .ZN(_0082_));
 INV_X1 _4631_ (.A(net90),
    .ZN(_0919_));
 NOR2_X1 _4632_ (.A1(rst),
    .A2(_0919_),
    .ZN(_0081_));
 NOR2_X1 _4633_ (.A1(rst),
    .A2(_1286_),
    .ZN(_0080_));
 AND2_X1 _4634_ (.A1(_1253_),
    .A2(net84),
    .ZN(_0079_));
 NOR2_X1 _4635_ (.A1(rst),
    .A2(_1550_),
    .ZN(_0078_));
 NOR2_X1 _4636_ (.A1(rst),
    .A2(_0330_),
    .ZN(_0077_));
 NOR2_X1 _4637_ (.A1(rst),
    .A2(_0749_),
    .ZN(_0076_));
 INV_X1 _4638_ (.A(net20),
    .ZN(_0920_));
 NOR2_X1 _4639_ (.A1(rst),
    .A2(net21),
    .ZN(_0075_));
 INV_X1 _4640_ (.A(net1),
    .ZN(_0921_));
 NOR2_X1 _4641_ (.A1(rst),
    .A2(net2),
    .ZN(_0074_));
 INV_X1 _4642_ (.A(net4),
    .ZN(_0922_));
 NOR2_X1 _4643_ (.A1(rst),
    .A2(net5),
    .ZN(_0073_));
 INV_X1 _4644_ (.A(net22),
    .ZN(_0923_));
 NOR2_X1 _4645_ (.A1(rst),
    .A2(net23),
    .ZN(_0072_));
 INV_X1 _4646_ (.A(net39),
    .ZN(_0924_));
 NOR2_X1 _4647_ (.A1(rst),
    .A2(net40),
    .ZN(_0071_));
 INV_X1 _4648_ (.A(net27),
    .ZN(_0925_));
 NOR2_X1 _4649_ (.A1(rst),
    .A2(net28),
    .ZN(_0070_));
 AND2_X1 _4650_ (.A1(_1253_),
    .A2(net25),
    .ZN(_0069_));
 INV_X1 _4651_ (.A(net7),
    .ZN(_0926_));
 NOR2_X1 _4652_ (.A1(rst),
    .A2(net8),
    .ZN(_0068_));
 AND2_X1 _4653_ (.A1(_1253_),
    .A2(net10),
    .ZN(_0067_));
 INV_X1 _4654_ (.A(net73),
    .ZN(_0927_));
 NOR2_X1 _4655_ (.A1(rst),
    .A2(net74),
    .ZN(_0066_));
 AND2_X1 _4656_ (.A1(_1253_),
    .A2(net12),
    .ZN(_0065_));
 INV_X1 _4657_ (.A(net33),
    .ZN(_0928_));
 NOR2_X1 _4658_ (.A1(rst),
    .A2(net34),
    .ZN(_0064_));
 INV_X1 _4659_ (.A(net35),
    .ZN(_0929_));
 NOR2_X1 _4660_ (.A1(rst),
    .A2(net36),
    .ZN(_0063_));
 INV_X1 _4661_ (.A(net43),
    .ZN(_0930_));
 NOR2_X1 _4662_ (.A1(rst),
    .A2(net44),
    .ZN(_0062_));
 INV_X1 _4663_ (.A(net37),
    .ZN(_0931_));
 NOR2_X1 _4664_ (.A1(rst),
    .A2(net38),
    .ZN(_0061_));
 INV_X1 _4665_ (.A(net17),
    .ZN(_0932_));
 NOR2_X1 _4666_ (.A1(rst),
    .A2(net18),
    .ZN(_0060_));
 INV_X1 _4667_ (.A(net14),
    .ZN(_0933_));
 NOR2_X1 _4668_ (.A1(rst),
    .A2(net15),
    .ZN(_0059_));
 INV_X1 _4669_ (.A(net31),
    .ZN(_0934_));
 NOR2_X1 _4670_ (.A1(rst),
    .A2(net32),
    .ZN(_0058_));
 INV_X1 _4671_ (.A(net47),
    .ZN(_0935_));
 NOR2_X1 _4672_ (.A1(rst),
    .A2(_0935_),
    .ZN(_0057_));
 INV_X1 _4673_ (.A(net45),
    .ZN(_0936_));
 NOR2_X1 _4674_ (.A1(rst),
    .A2(net46),
    .ZN(_0056_));
 AND2_X1 _4675_ (.A1(_1253_),
    .A2(net62),
    .ZN(_0055_));
 AND2_X1 _4676_ (.A1(_1253_),
    .A2(net29),
    .ZN(_0054_));
 AND2_X1 _4677_ (.A1(_1253_),
    .A2(x[9]),
    .ZN(_0053_));
 AND2_X1 _4678_ (.A1(_1253_),
    .A2(x[8]),
    .ZN(_0052_));
 AND2_X1 _4679_ (.A1(_1253_),
    .A2(x[7]),
    .ZN(_0051_));
 AND2_X1 _4680_ (.A1(_1253_),
    .A2(x[6]),
    .ZN(_0050_));
 AND2_X1 _4681_ (.A1(_1253_),
    .A2(x[5]),
    .ZN(_0049_));
 AND2_X1 _4682_ (.A1(_1253_),
    .A2(x[4]),
    .ZN(_0048_));
 AND2_X1 _4683_ (.A1(_1253_),
    .A2(x[3]),
    .ZN(_0047_));
 AND2_X1 _4684_ (.A1(_1253_),
    .A2(x[2]),
    .ZN(_0046_));
 AND2_X1 _4685_ (.A1(_1253_),
    .A2(x[1]),
    .ZN(_0045_));
 AND2_X1 _4686_ (.A1(_1253_),
    .A2(x[10]),
    .ZN(_0044_));
 AND2_X1 _4687_ (.A1(_1253_),
    .A2(x[0]),
    .ZN(_0043_));
 NAND2_X1 _4688_ (.A1(\section_1.yn2[9] ),
    .A2(\section_1.yn2[10] ),
    .ZN(_0937_));
 NAND2_X1 _4689_ (.A1(\section_1.yn2[8] ),
    .A2(\section_1.yn2[6] ),
    .ZN(_0938_));
 XOR2_X1 _4690_ (.A(\section_1.yn2[9] ),
    .B(\section_1.yn2[7] ),
    .Z(_0939_));
 XOR2_X1 _4691_ (.A(_0937_),
    .B(_0939_),
    .Z(_0940_));
 OAI22_X1 _4692_ (.A1(\section_1.yn2[7] ),
    .A2(_0937_),
    .B1(_0938_),
    .B2(_0940_),
    .ZN(_0941_));
 XOR2_X1 _4693_ (.A(\section_1.xn1[6] ),
    .B(\section_1.t1[1] ),
    .Z(_0942_));
 NAND3_X1 _4694_ (.A1(\section_1.xn1[5] ),
    .A2(\section_1.t1[0] ),
    .A3(_0942_),
    .ZN(_0943_));
 NAND2_X1 _4695_ (.A1(\section_1.xn1[6] ),
    .A2(\section_1.t1[1] ),
    .ZN(_0944_));
 XNOR2_X1 _4696_ (.A(\section_1.xn1[7] ),
    .B(\section_1.t1[2] ),
    .ZN(_0945_));
 XOR2_X1 _4697_ (.A(_0944_),
    .B(_0945_),
    .Z(_0946_));
 XNOR2_X1 _4698_ (.A(_0943_),
    .B(_0946_),
    .ZN(_0947_));
 XNOR2_X1 _4699_ (.A(\in_reg1[5] ),
    .B(_0947_),
    .ZN(_0948_));
 XNOR2_X1 _4700_ (.A(_0934_),
    .B(_0948_),
    .ZN(_0949_));
 NAND2_X1 _4701_ (.A1(\section_1.xn1[5] ),
    .A2(\section_1.t1[0] ),
    .ZN(_0950_));
 XNOR2_X1 _4702_ (.A(_0950_),
    .B(_0942_),
    .ZN(_0951_));
 XNOR2_X1 _4703_ (.A(\in_reg1[4] ),
    .B(_0951_),
    .ZN(_0952_));
 OR2_X1 _4704_ (.A1(_0935_),
    .A2(_0952_),
    .ZN(_0953_));
 NAND2_X1 _4705_ (.A1(\in_reg1[4] ),
    .A2(_0951_),
    .ZN(_0954_));
 AOI21_X1 _4706_ (.A(_0949_),
    .B1(_0953_),
    .B2(_0954_),
    .ZN(_0955_));
 AND3_X1 _4707_ (.A1(_0954_),
    .A2(_0953_),
    .A3(_0949_),
    .ZN(_0956_));
 OR2_X1 _4708_ (.A1(_0955_),
    .A2(_0956_),
    .ZN(_0957_));
 XNOR2_X1 _4709_ (.A(\in_reg1[3] ),
    .B(\section_1.xn2[5] ),
    .ZN(_0958_));
 NOR2_X1 _4710_ (.A1(_0957_),
    .A2(_0958_),
    .ZN(_0959_));
 NOR2_X1 _4711_ (.A1(_0955_),
    .A2(_0959_),
    .ZN(_0960_));
 OR2_X1 _4712_ (.A1(_0943_),
    .A2(_0945_),
    .ZN(_0961_));
 XNOR2_X1 _4713_ (.A(\section_1.xn1[8] ),
    .B(\section_1.t1[3] ),
    .ZN(_0962_));
 NAND2_X1 _4714_ (.A1(\section_1.xn1[7] ),
    .A2(\section_1.t1[2] ),
    .ZN(_0963_));
 OAI21_X1 _4715_ (.A(_0963_),
    .B1(_0945_),
    .B2(_0944_),
    .ZN(_0964_));
 XOR2_X1 _4716_ (.A(_0962_),
    .B(_0964_),
    .Z(_0965_));
 XNOR2_X1 _4717_ (.A(_0961_),
    .B(_0965_),
    .ZN(_0966_));
 XNOR2_X1 _4718_ (.A(_0931_),
    .B(_0966_),
    .ZN(_0967_));
 XNOR2_X1 _4719_ (.A(_0932_),
    .B(_0967_),
    .ZN(_0968_));
 OR2_X1 _4720_ (.A1(_0934_),
    .A2(_0948_),
    .ZN(_0969_));
 NAND2_X1 _4721_ (.A1(\in_reg1[5] ),
    .A2(_0947_),
    .ZN(_0970_));
 AOI21_X1 _4722_ (.A(_0968_),
    .B1(_0969_),
    .B2(_0970_),
    .ZN(_0971_));
 AND3_X1 _4723_ (.A1(_0970_),
    .A2(_0969_),
    .A3(_0968_),
    .ZN(_0972_));
 OR2_X1 _4724_ (.A1(_0971_),
    .A2(_0972_),
    .ZN(_0973_));
 XOR2_X1 _4725_ (.A(\in_reg1[4] ),
    .B(\section_1.xn2[6] ),
    .Z(_0974_));
 XNOR2_X1 _4726_ (.A(_0973_),
    .B(_0974_),
    .ZN(_0975_));
 XNOR2_X1 _4727_ (.A(_0960_),
    .B(_0975_),
    .ZN(_0976_));
 NAND2_X1 _4728_ (.A1(\section_1.xn2[3] ),
    .A2(\section_1.xn2[4] ),
    .ZN(_0977_));
 NAND2_X1 _4729_ (.A1(\in_reg1[3] ),
    .A2(\section_1.xn2[5] ),
    .ZN(_0978_));
 XOR2_X1 _4730_ (.A(\section_1.xn2[4] ),
    .B(\section_1.xn2[5] ),
    .Z(_0979_));
 XNOR2_X1 _4731_ (.A(_0978_),
    .B(_0979_),
    .ZN(_0980_));
 XNOR2_X1 _4732_ (.A(_0977_),
    .B(_0980_),
    .ZN(_0981_));
 XNOR2_X1 _4733_ (.A(_0976_),
    .B(_0981_),
    .ZN(_0982_));
 XNOR2_X1 _4734_ (.A(_0935_),
    .B(_0952_),
    .ZN(_0983_));
 XOR2_X1 _4735_ (.A(\section_1.xn1[5] ),
    .B(\section_1.t1[0] ),
    .Z(_0984_));
 XNOR2_X1 _4736_ (.A(\in_reg1[3] ),
    .B(_0984_),
    .ZN(_0985_));
 OR2_X1 _4737_ (.A1(_0936_),
    .A2(_0985_),
    .ZN(_0986_));
 NAND2_X1 _4738_ (.A1(\in_reg1[3] ),
    .A2(_0984_),
    .ZN(_0987_));
 AOI21_X1 _4739_ (.A(_0983_),
    .B1(_0986_),
    .B2(_0987_),
    .ZN(_0988_));
 AND3_X1 _4740_ (.A1(_0987_),
    .A2(_0986_),
    .A3(_0983_),
    .ZN(_0989_));
 OR2_X1 _4741_ (.A1(_0988_),
    .A2(_0989_),
    .ZN(_0990_));
 XNOR2_X1 _4742_ (.A(\in_reg1[2] ),
    .B(\section_1.xn2[4] ),
    .ZN(_0991_));
 NOR2_X1 _4743_ (.A1(_0990_),
    .A2(_0991_),
    .ZN(_0992_));
 NOR2_X1 _4744_ (.A1(_0988_),
    .A2(_0992_),
    .ZN(_0993_));
 XOR2_X1 _4745_ (.A(_0957_),
    .B(_0958_),
    .Z(_0994_));
 XNOR2_X1 _4746_ (.A(_0993_),
    .B(_0994_),
    .ZN(_0995_));
 NAND2_X1 _4747_ (.A1(\section_1.xn2[2] ),
    .A2(\section_1.xn2[3] ),
    .ZN(_0996_));
 NAND2_X1 _4748_ (.A1(\in_reg1[2] ),
    .A2(\section_1.xn2[4] ),
    .ZN(_0997_));
 XOR2_X1 _4749_ (.A(\section_1.xn2[3] ),
    .B(\section_1.xn2[4] ),
    .Z(_0998_));
 XNOR2_X1 _4750_ (.A(_0997_),
    .B(_0998_),
    .ZN(_0999_));
 XNOR2_X1 _4751_ (.A(_0996_),
    .B(_0999_),
    .ZN(_1000_));
 NAND2_X1 _4752_ (.A1(_0995_),
    .A2(_1000_),
    .ZN(_1001_));
 OAI21_X1 _4753_ (.A(_0994_),
    .B1(_0992_),
    .B2(_0988_),
    .ZN(_1002_));
 AOI21_X1 _4754_ (.A(_0982_),
    .B1(_1001_),
    .B2(_1002_),
    .ZN(_1003_));
 AND3_X1 _4755_ (.A1(_1002_),
    .A2(_1001_),
    .A3(_0982_),
    .ZN(_1004_));
 NOR2_X1 _4756_ (.A1(_1003_),
    .A2(_1004_),
    .ZN(_1005_));
 AOI21_X1 _4757_ (.A(_0998_),
    .B1(\section_1.xn2[4] ),
    .B2(\in_reg1[2] ),
    .ZN(_1006_));
 OAI22_X1 _4758_ (.A1(\section_1.xn2[3] ),
    .A2(_0997_),
    .B1(_0996_),
    .B2(_1006_),
    .ZN(_1007_));
 AOI21_X1 _4759_ (.A(_1003_),
    .B1(_1005_),
    .B2(_1007_),
    .ZN(_1008_));
 INV_X1 _4760_ (.A(_0973_),
    .ZN(_1009_));
 AOI21_X1 _4761_ (.A(_0971_),
    .B1(_1009_),
    .B2(_0974_),
    .ZN(_1010_));
 NOR2_X1 _4762_ (.A1(_0931_),
    .A2(_0966_),
    .ZN(_1011_));
 INV_X1 _4763_ (.A(_0967_),
    .ZN(_1012_));
 AOI21_X1 _4764_ (.A(_1011_),
    .B1(_1012_),
    .B2(\in_reg1[5] ),
    .ZN(_1013_));
 NOR2_X1 _4765_ (.A1(_0961_),
    .A2(_0965_),
    .ZN(_1014_));
 NOR3_X1 _4766_ (.A1(_0944_),
    .A2(_0945_),
    .A3(_0962_),
    .ZN(_1015_));
 XOR2_X1 _4767_ (.A(\section_1.xn1[9] ),
    .B(\section_1.t1[4] ),
    .Z(_1016_));
 NOR2_X1 _4768_ (.A1(_0963_),
    .A2(_0962_),
    .ZN(_1017_));
 AOI21_X1 _4769_ (.A(_1017_),
    .B1(\section_1.t1[3] ),
    .B2(\section_1.xn1[8] ),
    .ZN(_1018_));
 XNOR2_X1 _4770_ (.A(_1016_),
    .B(_1018_),
    .ZN(_1019_));
 XOR2_X1 _4771_ (.A(_1015_),
    .B(_1019_),
    .Z(_1020_));
 XNOR2_X1 _4772_ (.A(_1014_),
    .B(_1020_),
    .ZN(_1021_));
 XNOR2_X1 _4773_ (.A(_0930_),
    .B(_1021_),
    .ZN(_1022_));
 XNOR2_X1 _4774_ (.A(_0931_),
    .B(_1022_),
    .ZN(_1023_));
 XOR2_X1 _4775_ (.A(_1013_),
    .B(_1023_),
    .Z(_1024_));
 XOR2_X1 _4776_ (.A(\in_reg1[5] ),
    .B(\section_1.xn2[7] ),
    .Z(_1025_));
 XNOR2_X1 _4777_ (.A(_1024_),
    .B(_1025_),
    .ZN(_1026_));
 XOR2_X1 _4778_ (.A(_1010_),
    .B(_1026_),
    .Z(_1027_));
 AND2_X1 _4779_ (.A1(\section_1.xn2[4] ),
    .A2(\section_1.xn2[5] ),
    .ZN(_1028_));
 OR2_X1 _4780_ (.A1(\section_1.xn2[6] ),
    .A2(\section_1.xn2[5] ),
    .ZN(_1029_));
 NAND2_X1 _4781_ (.A1(\section_1.xn2[6] ),
    .A2(\section_1.xn2[5] ),
    .ZN(_1030_));
 AOI22_X1 _4782_ (.A1(\in_reg1[4] ),
    .A2(\section_1.xn2[6] ),
    .B1(_1029_),
    .B2(_1030_),
    .ZN(_1031_));
 INV_X1 _4783_ (.A(\section_1.xn2[6] ),
    .ZN(_1032_));
 NOR3_X1 _4784_ (.A1(_0934_),
    .A2(_1032_),
    .A3(\section_1.xn2[5] ),
    .ZN(_1033_));
 NOR2_X1 _4785_ (.A1(_1031_),
    .A2(_1033_),
    .ZN(_1034_));
 XOR2_X1 _4786_ (.A(_1028_),
    .B(_1034_),
    .Z(_1035_));
 XNOR2_X1 _4787_ (.A(_1027_),
    .B(_1035_),
    .ZN(_1036_));
 NAND2_X1 _4788_ (.A1(_0976_),
    .A2(_0981_),
    .ZN(_1037_));
 OAI21_X1 _4789_ (.A(_0975_),
    .B1(_0959_),
    .B2(_0955_),
    .ZN(_1038_));
 AOI21_X1 _4790_ (.A(_1036_),
    .B1(_1037_),
    .B2(_1038_),
    .ZN(_1039_));
 AND3_X1 _4791_ (.A1(_1038_),
    .A2(_1037_),
    .A3(_1036_),
    .ZN(_1040_));
 NOR2_X1 _4792_ (.A1(_1039_),
    .A2(_1040_),
    .ZN(_1041_));
 NAND3_X1 _4793_ (.A1(\section_1.xn2[3] ),
    .A2(\section_1.xn2[4] ),
    .A3(_0980_),
    .ZN(_1042_));
 OAI21_X1 _4794_ (.A(_1042_),
    .B1(_0978_),
    .B2(\section_1.xn2[4] ),
    .ZN(_1043_));
 XNOR2_X1 _4795_ (.A(_1041_),
    .B(_1043_),
    .ZN(_1044_));
 NOR2_X1 _4796_ (.A1(_1008_),
    .A2(_1044_),
    .ZN(_1045_));
 XOR2_X1 _4797_ (.A(_1008_),
    .B(_1044_),
    .Z(_1046_));
 NOR2_X1 _4798_ (.A1(_0925_),
    .A2(_0936_),
    .ZN(_1047_));
 XOR2_X1 _4799_ (.A(\section_1.t1[4] ),
    .B(\in_reg1[2] ),
    .Z(_1048_));
 AOI21_X1 _4800_ (.A(_1047_),
    .B1(_1048_),
    .B2(\in_reg1[1] ),
    .ZN(_1049_));
 XNOR2_X1 _4801_ (.A(_0936_),
    .B(_0985_),
    .ZN(_1050_));
 XOR2_X1 _4802_ (.A(_1049_),
    .B(_1050_),
    .Z(_1051_));
 XOR2_X1 _4803_ (.A(\in_reg1[1] ),
    .B(\section_1.xn2[3] ),
    .Z(_1052_));
 NAND2_X1 _4804_ (.A1(_1051_),
    .A2(_1052_),
    .ZN(_1053_));
 OAI21_X1 _4805_ (.A(_1053_),
    .B1(_1050_),
    .B2(_1049_),
    .ZN(_1054_));
 XOR2_X1 _4806_ (.A(_0990_),
    .B(_0991_),
    .Z(_1055_));
 XOR2_X1 _4807_ (.A(_1054_),
    .B(_1055_),
    .Z(_1056_));
 NAND2_X1 _4808_ (.A1(\section_1.xn2[1] ),
    .A2(\section_1.xn2[2] ),
    .ZN(_1057_));
 NAND2_X1 _4809_ (.A1(\in_reg1[1] ),
    .A2(\section_1.xn2[3] ),
    .ZN(_1058_));
 XOR2_X1 _4810_ (.A(\section_1.xn2[2] ),
    .B(\section_1.xn2[3] ),
    .Z(_1059_));
 XNOR2_X1 _4811_ (.A(_1058_),
    .B(_1059_),
    .ZN(_1060_));
 XNOR2_X1 _4812_ (.A(_1057_),
    .B(_1060_),
    .ZN(_1061_));
 AOI22_X1 _4813_ (.A1(_1054_),
    .A2(_1055_),
    .B1(_1056_),
    .B2(_1061_),
    .ZN(_1062_));
 XNOR2_X1 _4814_ (.A(_0995_),
    .B(_1000_),
    .ZN(_1063_));
 XOR2_X1 _4815_ (.A(_1062_),
    .B(_1063_),
    .Z(_1064_));
 AOI21_X1 _4816_ (.A(_1059_),
    .B1(\section_1.xn2[3] ),
    .B2(\in_reg1[1] ),
    .ZN(_1065_));
 OAI22_X1 _4817_ (.A1(\section_1.xn2[2] ),
    .A2(_1058_),
    .B1(_1057_),
    .B2(_1065_),
    .ZN(_1066_));
 NAND2_X1 _4818_ (.A1(_1064_),
    .A2(_1066_),
    .ZN(_1067_));
 OAI21_X1 _4819_ (.A(_1067_),
    .B1(_1063_),
    .B2(_1062_),
    .ZN(_1068_));
 XOR2_X1 _4820_ (.A(_1005_),
    .B(_1007_),
    .Z(_1069_));
 NAND2_X1 _4821_ (.A1(_1068_),
    .A2(_1069_),
    .ZN(_1070_));
 XOR2_X1 _4822_ (.A(_1064_),
    .B(_1066_),
    .Z(_1071_));
 XNOR2_X1 _4823_ (.A(\in_reg1[1] ),
    .B(_1048_),
    .ZN(_1072_));
 NOR2_X1 _4824_ (.A1(\section_1.t1[3] ),
    .A2(\in_reg1[1] ),
    .ZN(_1073_));
 AOI21_X1 _4825_ (.A(\in_reg1[0] ),
    .B1(\in_reg1[1] ),
    .B2(\section_1.t1[3] ),
    .ZN(_1074_));
 NOR3_X1 _4826_ (.A1(_1072_),
    .A2(_1073_),
    .A3(_1074_),
    .ZN(_1075_));
 NOR2_X1 _4827_ (.A1(_1073_),
    .A2(_1074_),
    .ZN(_1076_));
 XNOR2_X1 _4828_ (.A(_1072_),
    .B(_1076_),
    .ZN(_1077_));
 XOR2_X1 _4829_ (.A(\in_reg1[0] ),
    .B(\section_1.xn2[2] ),
    .Z(_1078_));
 AOI21_X1 _4830_ (.A(_1075_),
    .B1(_1077_),
    .B2(_1078_),
    .ZN(_1079_));
 XNOR2_X1 _4831_ (.A(_1051_),
    .B(_1052_),
    .ZN(_1080_));
 NOR2_X1 _4832_ (.A1(_1079_),
    .A2(_1080_),
    .ZN(_1081_));
 XOR2_X1 _4833_ (.A(_1079_),
    .B(_1080_),
    .Z(_1082_));
 NAND2_X1 _4834_ (.A1(\section_1.xn2[0] ),
    .A2(\section_1.xn2[1] ),
    .ZN(_1083_));
 NAND2_X1 _4835_ (.A1(\in_reg1[0] ),
    .A2(\section_1.xn2[2] ),
    .ZN(_1084_));
 XOR2_X1 _4836_ (.A(\section_1.xn2[1] ),
    .B(\section_1.xn2[2] ),
    .Z(_1085_));
 XNOR2_X1 _4837_ (.A(_1084_),
    .B(_1085_),
    .ZN(_1086_));
 XNOR2_X1 _4838_ (.A(_1083_),
    .B(_1086_),
    .ZN(_1087_));
 AOI21_X1 _4839_ (.A(_1081_),
    .B1(_1082_),
    .B2(_1087_),
    .ZN(_1088_));
 XNOR2_X1 _4840_ (.A(_1056_),
    .B(_1061_),
    .ZN(_1089_));
 XOR2_X1 _4841_ (.A(_1088_),
    .B(_1089_),
    .Z(_1090_));
 AOI21_X1 _4842_ (.A(_1085_),
    .B1(\section_1.xn2[2] ),
    .B2(\in_reg1[0] ),
    .ZN(_1091_));
 OAI22_X1 _4843_ (.A1(\section_1.xn2[1] ),
    .A2(_1084_),
    .B1(_1083_),
    .B2(_1091_),
    .ZN(_1092_));
 AND2_X1 _4844_ (.A1(_1090_),
    .A2(_1092_),
    .ZN(_1093_));
 NOR2_X1 _4845_ (.A1(_1088_),
    .A2(_1089_),
    .ZN(_1094_));
 OAI21_X1 _4846_ (.A(_1071_),
    .B1(_1093_),
    .B2(_1094_),
    .ZN(_1095_));
 INV_X1 _4847_ (.A(_1095_),
    .ZN(_1096_));
 NOR2_X1 _4848_ (.A1(_1094_),
    .A2(_1093_),
    .ZN(_1097_));
 XNOR2_X1 _4849_ (.A(_1097_),
    .B(_1071_),
    .ZN(_1098_));
 XOR2_X1 _4850_ (.A(_1090_),
    .B(_1092_),
    .Z(_1099_));
 INV_X1 _4851_ (.A(_1099_),
    .ZN(_1100_));
 INV_X1 _4852_ (.A(\section_1.xn2[0] ),
    .ZN(_1101_));
 XOR2_X1 _4853_ (.A(\section_1.t1[2] ),
    .B(\in_reg1[0] ),
    .Z(_1102_));
 NAND2_X1 _4854_ (.A1(\section_1.xn2[0] ),
    .A2(_1102_),
    .ZN(_1103_));
 XOR2_X1 _4855_ (.A(\section_1.t1[3] ),
    .B(\in_reg1[1] ),
    .Z(_1104_));
 NAND2_X1 _4856_ (.A1(_0926_),
    .A2(\in_reg1[0] ),
    .ZN(_1105_));
 XNOR2_X1 _4857_ (.A(_1104_),
    .B(_1105_),
    .ZN(_1106_));
 XNOR2_X1 _4858_ (.A(\section_1.xn2[1] ),
    .B(_1106_),
    .ZN(_1107_));
 AOI21_X1 _4859_ (.A(_1101_),
    .B1(_1103_),
    .B2(_1107_),
    .ZN(_1108_));
 NAND2_X1 _4860_ (.A1(\section_1.xn2[1] ),
    .A2(_1106_),
    .ZN(_1109_));
 NAND2_X1 _4861_ (.A1(\section_1.t1[2] ),
    .A2(\in_reg1[0] ),
    .ZN(_1110_));
 OAI21_X1 _4862_ (.A(_1109_),
    .B1(_1110_),
    .B2(_1104_),
    .ZN(_1111_));
 XNOR2_X1 _4863_ (.A(_1077_),
    .B(_1078_),
    .ZN(_1112_));
 INV_X1 _4864_ (.A(_1112_),
    .ZN(_1113_));
 XNOR2_X1 _4865_ (.A(_1111_),
    .B(_1113_),
    .ZN(_1114_));
 XNOR2_X1 _4866_ (.A(\section_1.xn2[0] ),
    .B(\section_1.xn2[1] ),
    .ZN(_1115_));
 XOR2_X1 _4867_ (.A(_1114_),
    .B(_1115_),
    .Z(_1116_));
 AND2_X1 _4868_ (.A1(_1108_),
    .A2(_1116_),
    .ZN(_1117_));
 XNOR2_X1 _4869_ (.A(_1082_),
    .B(_1087_),
    .ZN(_1118_));
 OR2_X1 _4870_ (.A1(_1114_),
    .A2(_1115_),
    .ZN(_1119_));
 NAND2_X1 _4871_ (.A1(_1111_),
    .A2(_1113_),
    .ZN(_1120_));
 AOI21_X1 _4872_ (.A(_1118_),
    .B1(_1119_),
    .B2(_1120_),
    .ZN(_1121_));
 INV_X1 _4873_ (.A(_1121_),
    .ZN(_1122_));
 NAND3_X1 _4874_ (.A1(_1120_),
    .A2(_1119_),
    .A3(_1118_),
    .ZN(_1123_));
 AND2_X1 _4875_ (.A1(_1122_),
    .A2(_1123_),
    .ZN(_1124_));
 NAND2_X1 _4876_ (.A1(_1117_),
    .A2(_1124_),
    .ZN(_1125_));
 AOI21_X1 _4877_ (.A(_1100_),
    .B1(_1125_),
    .B2(_1122_),
    .ZN(_1126_));
 AOI21_X1 _4878_ (.A(_1096_),
    .B1(_1098_),
    .B2(_1126_),
    .ZN(_1127_));
 XNOR2_X1 _4879_ (.A(_1068_),
    .B(_1069_),
    .ZN(_1128_));
 OAI21_X1 _4880_ (.A(_1070_),
    .B1(_1127_),
    .B2(_1128_),
    .ZN(_1129_));
 AOI21_X1 _4881_ (.A(_1045_),
    .B1(_1046_),
    .B2(_1129_),
    .ZN(_1130_));
 AOI21_X1 _4882_ (.A(_1039_),
    .B1(_1041_),
    .B2(_1043_),
    .ZN(_1131_));
 AOI21_X1 _4883_ (.A(_1033_),
    .B1(_1034_),
    .B2(_1028_),
    .ZN(_1132_));
 NOR2_X1 _4884_ (.A1(_1010_),
    .A2(_1026_),
    .ZN(_1133_));
 AOI21_X1 _4885_ (.A(_1133_),
    .B1(_1027_),
    .B2(_1035_),
    .ZN(_1134_));
 NAND2_X1 _4886_ (.A1(\in_reg1[5] ),
    .A2(\section_1.xn2[7] ),
    .ZN(_1135_));
 XOR2_X1 _4887_ (.A(\section_1.xn2[7] ),
    .B(\section_1.xn2[6] ),
    .Z(_1136_));
 XNOR2_X1 _4888_ (.A(_1135_),
    .B(_1136_),
    .ZN(_1137_));
 XNOR2_X1 _4889_ (.A(_1030_),
    .B(_1137_),
    .ZN(_1138_));
 NOR2_X1 _4890_ (.A1(_1013_),
    .A2(_1023_),
    .ZN(_1139_));
 AOI21_X1 _4891_ (.A(_1139_),
    .B1(_1024_),
    .B2(_1025_),
    .ZN(_1140_));
 XOR2_X1 _4892_ (.A(\in_reg1[6] ),
    .B(\section_1.xn2[8] ),
    .Z(_1141_));
 NOR2_X1 _4893_ (.A1(_0930_),
    .A2(_1021_),
    .ZN(_1142_));
 INV_X1 _4894_ (.A(_1022_),
    .ZN(_1143_));
 AOI21_X1 _4895_ (.A(_1142_),
    .B1(_1143_),
    .B2(\in_reg1[6] ),
    .ZN(_1144_));
 NAND2_X1 _4896_ (.A1(_1015_),
    .A2(_1019_),
    .ZN(_1145_));
 NAND2_X1 _4897_ (.A1(_1014_),
    .A2(_1020_),
    .ZN(_1146_));
 NAND2_X1 _4898_ (.A1(_1145_),
    .A2(_1146_),
    .ZN(_1147_));
 NAND2_X1 _4899_ (.A1(_1017_),
    .A2(_1016_),
    .ZN(_1148_));
 XOR2_X1 _4900_ (.A(\section_1.xn1[5] ),
    .B(\section_1.xn1[10] ),
    .Z(_1149_));
 NAND3_X1 _4901_ (.A1(\section_1.xn1[8] ),
    .A2(\section_1.t1[3] ),
    .A3(_1016_),
    .ZN(_1150_));
 OAI21_X1 _4902_ (.A(_1150_),
    .B1(_0925_),
    .B2(_0920_),
    .ZN(_1151_));
 XOR2_X1 _4903_ (.A(_1149_),
    .B(_1151_),
    .Z(_1152_));
 XOR2_X1 _4904_ (.A(_1148_),
    .B(_1152_),
    .Z(_1153_));
 XNOR2_X1 _4905_ (.A(_1147_),
    .B(_1153_),
    .ZN(_1154_));
 XNOR2_X1 _4906_ (.A(\in_reg1[8] ),
    .B(_1154_),
    .ZN(_1155_));
 XNOR2_X1 _4907_ (.A(_0930_),
    .B(_1155_),
    .ZN(_1156_));
 XOR2_X1 _4908_ (.A(_1144_),
    .B(_1156_),
    .Z(_1157_));
 XNOR2_X1 _4909_ (.A(_1141_),
    .B(_1157_),
    .ZN(_1158_));
 XOR2_X1 _4910_ (.A(_1140_),
    .B(_1158_),
    .Z(_1159_));
 XNOR2_X1 _4911_ (.A(_1138_),
    .B(_1159_),
    .ZN(_1160_));
 XNOR2_X1 _4912_ (.A(_1134_),
    .B(_1160_),
    .ZN(_1161_));
 XNOR2_X1 _4913_ (.A(_1132_),
    .B(_1161_),
    .ZN(_1162_));
 XNOR2_X1 _4914_ (.A(_1131_),
    .B(_1162_),
    .ZN(_1163_));
 XOR2_X1 _4915_ (.A(_1130_),
    .B(_1163_),
    .Z(_1164_));
 XNOR2_X1 _4916_ (.A(_0330_),
    .B(_1164_),
    .ZN(_1165_));
 NAND2_X1 _4917_ (.A1(\coll_reg[0] ),
    .A2(_1165_),
    .ZN(_1166_));
 INV_X1 _4918_ (.A(_1164_),
    .ZN(_1167_));
 OAI21_X1 _4919_ (.A(_1166_),
    .B1(_1167_),
    .B2(_0006_),
    .ZN(_1168_));
 OAI22_X1 _4920_ (.A1(_1134_),
    .A2(_1160_),
    .B1(_1161_),
    .B2(_1132_),
    .ZN(_1169_));
 NAND3_X1 _4921_ (.A1(\section_1.xn2[6] ),
    .A2(\section_1.xn2[5] ),
    .A3(_1137_),
    .ZN(_1170_));
 OAI21_X1 _4922_ (.A(_1170_),
    .B1(_1135_),
    .B2(\section_1.xn2[6] ),
    .ZN(_1171_));
 NOR2_X1 _4923_ (.A1(_1140_),
    .A2(_1158_),
    .ZN(_1172_));
 AOI21_X1 _4924_ (.A(_1172_),
    .B1(_1159_),
    .B2(_1138_),
    .ZN(_1173_));
 INV_X1 _4925_ (.A(_1173_),
    .ZN(_1174_));
 INV_X1 _4926_ (.A(\section_1.xn2[8] ),
    .ZN(_1175_));
 OAI211_X1 _4927_ (.A(\section_1.xn2[7] ),
    .B(\section_1.xn2[6] ),
    .C1(\in_reg1[6] ),
    .C2(_1175_),
    .ZN(_1176_));
 NAND2_X1 _4928_ (.A1(\in_reg1[6] ),
    .A2(\section_1.xn2[8] ),
    .ZN(_1177_));
 XNOR2_X1 _4929_ (.A(\section_1.xn2[8] ),
    .B(\section_1.xn2[7] ),
    .ZN(_1178_));
 XNOR2_X1 _4930_ (.A(_1177_),
    .B(_1178_),
    .ZN(_1179_));
 INV_X1 _4931_ (.A(\section_1.xn2[7] ),
    .ZN(_1180_));
 OAI21_X1 _4932_ (.A(_1179_),
    .B1(_1032_),
    .B2(_1180_),
    .ZN(_1181_));
 AND2_X1 _4933_ (.A1(_1176_),
    .A2(_1181_),
    .ZN(_1182_));
 NOR2_X1 _4934_ (.A1(_1144_),
    .A2(_1156_),
    .ZN(_1183_));
 AOI21_X1 _4935_ (.A(_1183_),
    .B1(_1157_),
    .B2(_1141_),
    .ZN(_1184_));
 XOR2_X1 _4936_ (.A(\in_reg1[7] ),
    .B(\section_1.xn2[9] ),
    .Z(_1185_));
 NOR2_X1 _4937_ (.A1(_0930_),
    .A2(_1155_),
    .ZN(_1186_));
 AOI21_X1 _4938_ (.A(_1186_),
    .B1(_1154_),
    .B2(\in_reg1[8] ),
    .ZN(_1187_));
 INV_X1 _4939_ (.A(_1150_),
    .ZN(_1188_));
 NAND2_X1 _4940_ (.A1(_1188_),
    .A2(_1149_),
    .ZN(_1189_));
 NAND3_X1 _4941_ (.A1(\section_1.xn1[9] ),
    .A2(\section_1.t1[4] ),
    .A3(_1149_),
    .ZN(_1190_));
 NOR3_X1 _4942_ (.A1(\section_1.xn1[6] ),
    .A2(_0924_),
    .A3(_0927_),
    .ZN(_1191_));
 NAND2_X1 _4943_ (.A1(_0923_),
    .A2(\section_1.xn1[10] ),
    .ZN(_1192_));
 MUX2_X1 _4944_ (.A(_0923_),
    .B(_0924_),
    .S(\section_1.xn1[10] ),
    .Z(_1193_));
 AOI21_X1 _4945_ (.A(_1191_),
    .B1(_1192_),
    .B2(_1193_),
    .ZN(_1194_));
 XNOR2_X1 _4946_ (.A(_1190_),
    .B(_1194_),
    .ZN(_1195_));
 XNOR2_X1 _4947_ (.A(_1189_),
    .B(_1195_),
    .ZN(_1196_));
 AOI21_X1 _4948_ (.A(_1153_),
    .B1(_1146_),
    .B2(_1145_),
    .ZN(_1197_));
 AND3_X1 _4949_ (.A1(_1017_),
    .A2(_1016_),
    .A3(_1152_),
    .ZN(_1198_));
 OAI21_X1 _4950_ (.A(_1196_),
    .B1(_1197_),
    .B2(_1198_),
    .ZN(_1199_));
 OR3_X1 _4951_ (.A1(_1198_),
    .A2(_1197_),
    .A3(_1196_),
    .ZN(_1200_));
 AND2_X1 _4952_ (.A1(_1199_),
    .A2(_1200_),
    .ZN(_1201_));
 XNOR2_X1 _4953_ (.A(\in_reg1[9] ),
    .B(_1201_),
    .ZN(_1202_));
 XNOR2_X1 _4954_ (.A(_0929_),
    .B(_1202_),
    .ZN(_1203_));
 XOR2_X1 _4955_ (.A(_1187_),
    .B(_1203_),
    .Z(_1204_));
 XNOR2_X1 _4956_ (.A(_1185_),
    .B(_1204_),
    .ZN(_1205_));
 XOR2_X1 _4957_ (.A(_1184_),
    .B(_1205_),
    .Z(_1206_));
 XOR2_X1 _4958_ (.A(_1182_),
    .B(_1206_),
    .Z(_1207_));
 XNOR2_X1 _4959_ (.A(_1174_),
    .B(_1207_),
    .ZN(_1208_));
 XNOR2_X1 _4960_ (.A(_1171_),
    .B(_1208_),
    .ZN(_1209_));
 NAND2_X1 _4961_ (.A1(_1169_),
    .A2(_1209_),
    .ZN(_1210_));
 OR2_X1 _4962_ (.A1(_1169_),
    .A2(_1209_),
    .ZN(_1211_));
 NAND2_X1 _4963_ (.A1(_1210_),
    .A2(_1211_),
    .ZN(_1212_));
 NOR2_X1 _4964_ (.A1(_1131_),
    .A2(_1162_),
    .ZN(_1213_));
 NOR2_X1 _4965_ (.A1(_1130_),
    .A2(_1163_),
    .ZN(_1214_));
 NOR2_X1 _4966_ (.A1(_1213_),
    .A2(_1214_),
    .ZN(_1215_));
 XNOR2_X1 _4967_ (.A(_1212_),
    .B(_1215_),
    .ZN(_1216_));
 XNOR2_X1 _4968_ (.A(\coll_reg[1] ),
    .B(_1216_),
    .ZN(_1217_));
 NAND2_X1 _4969_ (.A1(_1168_),
    .A2(_1217_),
    .ZN(_1218_));
 XOR2_X1 _4970_ (.A(_1168_),
    .B(_1217_),
    .Z(_1219_));
 NAND2_X1 _4971_ (.A1(\coll_reg[2] ),
    .A2(_1219_),
    .ZN(_1220_));
 NAND2_X1 _4972_ (.A1(_1218_),
    .A2(_1220_),
    .ZN(_1221_));
 NAND2_X1 _4973_ (.A1(_1561_),
    .A2(_1660_),
    .ZN(_1222_));
 OR2_X1 _4974_ (.A1(_1550_),
    .A2(_1216_),
    .ZN(_1223_));
 NAND3_X1 _4975_ (.A1(_1214_),
    .A2(_1210_),
    .A3(_1211_),
    .ZN(_1224_));
 INV_X1 _4976_ (.A(_1210_),
    .ZN(_1225_));
 AOI21_X1 _4977_ (.A(_1225_),
    .B1(_1211_),
    .B2(_1213_),
    .ZN(_1226_));
 INV_X1 _4978_ (.A(_1171_),
    .ZN(_1227_));
 NOR2_X1 _4979_ (.A1(_1227_),
    .A2(_1208_),
    .ZN(_1228_));
 AOI21_X1 _4980_ (.A(_1228_),
    .B1(_1207_),
    .B2(_1174_),
    .ZN(_1229_));
 OAI21_X1 _4981_ (.A(_1176_),
    .B1(_1177_),
    .B2(\section_1.xn2[7] ),
    .ZN(_1230_));
 INV_X1 _4982_ (.A(_1230_),
    .ZN(_1231_));
 NOR2_X1 _4983_ (.A1(_1184_),
    .A2(_1205_),
    .ZN(_1232_));
 AOI21_X1 _4984_ (.A(_1232_),
    .B1(_1206_),
    .B2(_1182_),
    .ZN(_1233_));
 INV_X1 _4985_ (.A(\section_1.xn2[9] ),
    .ZN(_1234_));
 OAI211_X1 _4986_ (.A(\section_1.xn2[8] ),
    .B(\section_1.xn2[7] ),
    .C1(\in_reg1[7] ),
    .C2(_1234_),
    .ZN(_1235_));
 NAND2_X1 _4987_ (.A1(\in_reg1[7] ),
    .A2(\section_1.xn2[9] ),
    .ZN(_1236_));
 XNOR2_X1 _4988_ (.A(\section_1.xn2[9] ),
    .B(\section_1.xn2[8] ),
    .ZN(_1237_));
 XNOR2_X1 _4989_ (.A(_1236_),
    .B(_1237_),
    .ZN(_1238_));
 OAI21_X1 _4990_ (.A(_1238_),
    .B1(_1180_),
    .B2(_1175_),
    .ZN(_1239_));
 AND2_X1 _4991_ (.A1(_1235_),
    .A2(_1239_),
    .ZN(_1240_));
 NOR2_X1 _4992_ (.A1(_1187_),
    .A2(_1203_),
    .ZN(_1241_));
 AOI21_X1 _4993_ (.A(_1241_),
    .B1(_1204_),
    .B2(_1185_),
    .ZN(_1242_));
 XOR2_X1 _4994_ (.A(\in_reg1[8] ),
    .B(\section_1.xn2[10] ),
    .Z(_1243_));
 INV_X1 _4995_ (.A(_1243_),
    .ZN(_1244_));
 NAND2_X1 _4996_ (.A1(\in_reg1[9] ),
    .A2(_1201_),
    .ZN(_1245_));
 OAI21_X1 _4997_ (.A(_1245_),
    .B1(_1202_),
    .B2(_0929_),
    .ZN(_1246_));
 INV_X1 _4998_ (.A(_1246_),
    .ZN(_1247_));
 NAND3_X1 _4999_ (.A1(_1188_),
    .A2(_1149_),
    .A3(_1195_),
    .ZN(_1248_));
 AOI211_X1 _5000_ (.A(_1190_),
    .B(_1191_),
    .C1(_1192_),
    .C2(_1193_),
    .ZN(_1249_));
 NAND4_X1 _5001_ (.A1(_0922_),
    .A2(_0923_),
    .A3(_0924_),
    .A4(\section_1.xn1[10] ),
    .ZN(_1250_));
 OAI21_X1 _5002_ (.A(\section_1.xn1[7] ),
    .B1(\section_1.xn1[5] ),
    .B2(_1192_),
    .ZN(_1251_));
 AND2_X1 _5003_ (.A1(_1250_),
    .A2(_1251_),
    .ZN(_1252_));
 XOR2_X1 _5004_ (.A(_1249_),
    .B(_1252_),
    .Z(_1254_));
 AND3_X1 _5005_ (.A1(_1248_),
    .A2(_1199_),
    .A3(_1254_),
    .ZN(_1255_));
 AOI21_X1 _5006_ (.A(_1254_),
    .B1(_1199_),
    .B2(_1248_),
    .ZN(_1256_));
 OR2_X1 _5007_ (.A1(_1255_),
    .A2(_1256_),
    .ZN(_1257_));
 XNOR2_X1 _5008_ (.A(_0933_),
    .B(_1257_),
    .ZN(_1258_));
 XNOR2_X1 _5009_ (.A(_0928_),
    .B(_1258_),
    .ZN(_1259_));
 XNOR2_X1 _5010_ (.A(_1247_),
    .B(_1259_),
    .ZN(_1260_));
 XNOR2_X1 _5011_ (.A(_1244_),
    .B(_1260_),
    .ZN(_1261_));
 XOR2_X1 _5012_ (.A(_1242_),
    .B(_1261_),
    .Z(_1262_));
 XNOR2_X1 _5013_ (.A(_1240_),
    .B(_1262_),
    .ZN(_1263_));
 XNOR2_X1 _5014_ (.A(_1233_),
    .B(_1263_),
    .ZN(_1265_));
 XNOR2_X1 _5015_ (.A(_1231_),
    .B(_1265_),
    .ZN(_1266_));
 XNOR2_X1 _5016_ (.A(_1229_),
    .B(_1266_),
    .ZN(_1267_));
 AND3_X1 _5017_ (.A1(_1224_),
    .A2(_1226_),
    .A3(_1267_),
    .ZN(_1268_));
 AOI21_X1 _5018_ (.A(_1267_),
    .B1(_1226_),
    .B2(_1224_),
    .ZN(_1269_));
 OR2_X1 _5019_ (.A1(_1268_),
    .A2(_1269_),
    .ZN(_1270_));
 XOR2_X1 _5020_ (.A(_1223_),
    .B(_1270_),
    .Z(_1271_));
 XNOR2_X1 _5021_ (.A(_1222_),
    .B(_1271_),
    .ZN(_1272_));
 AND2_X1 _5022_ (.A1(_1221_),
    .A2(_1272_),
    .ZN(_1273_));
 XOR2_X1 _5023_ (.A(_1221_),
    .B(_1272_),
    .Z(_1274_));
 AND2_X1 _5024_ (.A1(\coll_reg[7] ),
    .A2(_1274_),
    .ZN(_1276_));
 NOR2_X1 _5025_ (.A1(_1273_),
    .A2(_1276_),
    .ZN(_1277_));
 NAND3_X1 _5026_ (.A1(_1561_),
    .A2(_1660_),
    .A3(_1271_),
    .ZN(_1278_));
 OAI21_X1 _5027_ (.A(_1278_),
    .B1(_1270_),
    .B2(_1223_),
    .ZN(_1279_));
 NOR2_X1 _5028_ (.A1(_1229_),
    .A2(_1266_),
    .ZN(_1280_));
 NOR2_X1 _5029_ (.A1(_1280_),
    .A2(_1269_),
    .ZN(_1281_));
 OAI21_X1 _5030_ (.A(_1235_),
    .B1(_1236_),
    .B2(\section_1.xn2[8] ),
    .ZN(_1282_));
 NOR2_X1 _5031_ (.A1(_1242_),
    .A2(_1261_),
    .ZN(_1283_));
 AOI21_X1 _5032_ (.A(_1283_),
    .B1(_1262_),
    .B2(_1240_),
    .ZN(_1284_));
 INV_X1 _5033_ (.A(\section_1.xn2[10] ),
    .ZN(_1285_));
 OAI211_X1 _5034_ (.A(\section_1.xn2[9] ),
    .B(\section_1.xn2[8] ),
    .C1(\in_reg1[8] ),
    .C2(_1285_),
    .ZN(_1287_));
 NAND2_X1 _5035_ (.A1(\in_reg1[8] ),
    .A2(\section_1.xn2[10] ),
    .ZN(_1288_));
 XNOR2_X1 _5036_ (.A(\section_1.xn2[10] ),
    .B(\section_1.xn2[9] ),
    .ZN(_1289_));
 XNOR2_X1 _5037_ (.A(_1288_),
    .B(_1289_),
    .ZN(_1290_));
 OAI21_X1 _5038_ (.A(_1290_),
    .B1(_1175_),
    .B2(_1234_),
    .ZN(_1291_));
 AND2_X1 _5039_ (.A1(_1287_),
    .A2(_1291_),
    .ZN(_1292_));
 OR2_X1 _5040_ (.A1(_1247_),
    .A2(_1259_),
    .ZN(_1293_));
 OAI21_X1 _5041_ (.A(_1293_),
    .B1(_1260_),
    .B2(_1244_),
    .ZN(_1294_));
 NOR2_X1 _5042_ (.A1(\in_reg1[9] ),
    .A2(\section_1.xn2[10] ),
    .ZN(_1295_));
 NOR2_X1 _5043_ (.A1(_0928_),
    .A2(_1285_),
    .ZN(_1296_));
 NOR2_X1 _5044_ (.A1(_1295_),
    .A2(_1296_),
    .ZN(_1298_));
 OAI22_X1 _5045_ (.A1(_0010_),
    .A2(_1257_),
    .B1(_1258_),
    .B2(_0928_),
    .ZN(_1299_));
 NOR3_X1 _5046_ (.A1(\section_1.xn1[8] ),
    .A2(\section_1.xn1[7] ),
    .A3(_1192_),
    .ZN(_1300_));
 AND2_X1 _5047_ (.A1(\section_1.xn1[5] ),
    .A2(_1300_),
    .ZN(_1301_));
 AOI21_X1 _5048_ (.A(_1300_),
    .B1(_1250_),
    .B2(\section_1.xn1[8] ),
    .ZN(_1302_));
 NOR2_X1 _5049_ (.A1(_1301_),
    .A2(_1302_),
    .ZN(_1303_));
 INV_X1 _5050_ (.A(_1252_),
    .ZN(_1304_));
 AOI21_X1 _5051_ (.A(_1256_),
    .B1(_1304_),
    .B2(_1249_),
    .ZN(_1305_));
 XNOR2_X1 _5052_ (.A(_1303_),
    .B(_1305_),
    .ZN(_1306_));
 XNOR2_X1 _5053_ (.A(_1299_),
    .B(_1306_),
    .ZN(_1307_));
 XNOR2_X1 _5054_ (.A(_1298_),
    .B(_1307_),
    .ZN(_1309_));
 XOR2_X1 _5055_ (.A(_1294_),
    .B(_1309_),
    .Z(_1310_));
 XNOR2_X1 _5056_ (.A(_1292_),
    .B(_1310_),
    .ZN(_1311_));
 XNOR2_X1 _5057_ (.A(_1284_),
    .B(_1311_),
    .ZN(_1312_));
 XNOR2_X1 _5058_ (.A(_1282_),
    .B(_1312_),
    .ZN(_1313_));
 NOR2_X1 _5059_ (.A1(_1231_),
    .A2(_1265_),
    .ZN(_1314_));
 OR2_X1 _5060_ (.A1(_1233_),
    .A2(_1263_),
    .ZN(_1315_));
 INV_X1 _5061_ (.A(_1315_),
    .ZN(_1316_));
 OAI21_X1 _5062_ (.A(_1313_),
    .B1(_1314_),
    .B2(_1316_),
    .ZN(_1317_));
 OR3_X1 _5063_ (.A1(_1316_),
    .A2(_1314_),
    .A3(_1313_),
    .ZN(_1318_));
 NAND2_X1 _5064_ (.A1(_1317_),
    .A2(_1318_),
    .ZN(_1320_));
 XOR2_X1 _5065_ (.A(_1281_),
    .B(_1320_),
    .Z(_1321_));
 XOR2_X1 _5066_ (.A(_1594_),
    .B(_1321_),
    .Z(_1322_));
 XNOR2_X1 _5067_ (.A(_1279_),
    .B(_1322_),
    .ZN(_1323_));
 XOR2_X1 _5068_ (.A(_1561_),
    .B(_1323_),
    .Z(_1324_));
 XOR2_X1 _5069_ (.A(_1277_),
    .B(_1324_),
    .Z(_1325_));
 XOR2_X1 _5070_ (.A(_0005_),
    .B(_2733_),
    .Z(_1326_));
 XNOR2_X1 _5071_ (.A(_1325_),
    .B(_1326_),
    .ZN(_1327_));
 NAND2_X1 _5072_ (.A1(\coll_reg[10] ),
    .A2(_2513_),
    .ZN(_1328_));
 XNOR2_X1 _5073_ (.A(\coll_reg[2] ),
    .B(_1219_),
    .ZN(_1329_));
 XOR2_X1 _5074_ (.A(_1129_),
    .B(_1046_),
    .Z(_1331_));
 NOR2_X1 _5075_ (.A1(_0749_),
    .A2(_1331_),
    .ZN(_1332_));
 XOR2_X1 _5076_ (.A(_1165_),
    .B(_1332_),
    .Z(_1333_));
 NAND2_X1 _5077_ (.A1(\coll_reg[1] ),
    .A2(_1333_),
    .ZN(_1334_));
 NAND2_X1 _5078_ (.A1(\coll_reg[0] ),
    .A2(_1331_),
    .ZN(_1335_));
 OR2_X1 _5079_ (.A1(_1335_),
    .A2(_1165_),
    .ZN(_1336_));
 AOI21_X1 _5080_ (.A(_1329_),
    .B1(_1334_),
    .B2(_1336_),
    .ZN(_1337_));
 NAND2_X1 _5081_ (.A1(_1336_),
    .A2(_1334_),
    .ZN(_1338_));
 XNOR2_X1 _5082_ (.A(_1338_),
    .B(_1329_),
    .ZN(_1339_));
 AND2_X1 _5083_ (.A1(\coll_reg[6] ),
    .A2(_1339_),
    .ZN(_1340_));
 NOR2_X1 _5084_ (.A1(_1337_),
    .A2(_1340_),
    .ZN(_1342_));
 XNOR2_X1 _5085_ (.A(_0918_),
    .B(_1274_),
    .ZN(_1343_));
 XNOR2_X1 _5086_ (.A(_1342_),
    .B(_1343_),
    .ZN(_1344_));
 OAI211_X1 _5087_ (.A(_1328_),
    .B(_1344_),
    .C1(\coll_reg[9] ),
    .C2(\coll_reg[10] ),
    .ZN(_1345_));
 OAI21_X1 _5088_ (.A(_1343_),
    .B1(_1340_),
    .B2(_1337_),
    .ZN(_1346_));
 AOI21_X1 _5089_ (.A(_1327_),
    .B1(_1345_),
    .B2(_1346_),
    .ZN(_1347_));
 NOR3_X1 _5090_ (.A1(\coll_reg[9] ),
    .A2(_0005_),
    .A3(_2732_),
    .ZN(_1348_));
 OAI21_X1 _5091_ (.A(_1324_),
    .B1(_1276_),
    .B2(_1273_),
    .ZN(_1349_));
 OR2_X1 _5092_ (.A1(_1325_),
    .A2(_1326_),
    .ZN(_1350_));
 NAND2_X1 _5093_ (.A1(_1349_),
    .A2(_1350_),
    .ZN(_1351_));
 XNOR2_X1 _5094_ (.A(\coll_reg[5] ),
    .B(_1924_),
    .ZN(_1353_));
 AND2_X1 _5095_ (.A1(_1594_),
    .A2(_1321_),
    .ZN(_1354_));
 OAI21_X1 _5096_ (.A(_1317_),
    .B1(_1320_),
    .B2(_1281_),
    .ZN(_1355_));
 OAI21_X1 _5097_ (.A(_1287_),
    .B1(_1288_),
    .B2(\section_1.xn2[9] ),
    .ZN(_1356_));
 AOI22_X1 _5098_ (.A1(_1294_),
    .A2(_1309_),
    .B1(_1310_),
    .B2(_1292_),
    .ZN(_1357_));
 OAI21_X1 _5099_ (.A(\section_1.xn2[10] ),
    .B1(\section_1.xn2[9] ),
    .B2(\in_reg1[9] ),
    .ZN(_1358_));
 AOI21_X1 _5100_ (.A(_1358_),
    .B1(_1296_),
    .B2(\section_1.xn2[9] ),
    .ZN(_1359_));
 NOR3_X1 _5101_ (.A1(_1295_),
    .A2(_1296_),
    .A3(_1307_),
    .ZN(_1360_));
 AOI21_X1 _5102_ (.A(_1360_),
    .B1(_1306_),
    .B2(_1299_),
    .ZN(_1361_));
 XOR2_X1 _5103_ (.A(\in_reg1[10] ),
    .B(\section_1.xn2[10] ),
    .Z(_1362_));
 INV_X1 _5104_ (.A(_0010_),
    .ZN(_1364_));
 NOR2_X1 _5105_ (.A1(_1302_),
    .A2(_1305_),
    .ZN(_1365_));
 XNOR2_X1 _5106_ (.A(_0920_),
    .B(_1300_),
    .ZN(_1366_));
 OR3_X1 _5107_ (.A1(_1301_),
    .A2(_1365_),
    .A3(_1366_),
    .ZN(_1367_));
 OAI21_X1 _5108_ (.A(_1366_),
    .B1(_1365_),
    .B2(_1301_),
    .ZN(_1368_));
 NAND2_X1 _5109_ (.A1(_1367_),
    .A2(_1368_),
    .ZN(_1369_));
 XNOR2_X1 _5110_ (.A(_1364_),
    .B(_1369_),
    .ZN(_1370_));
 XNOR2_X1 _5111_ (.A(_1362_),
    .B(_1370_),
    .ZN(_1371_));
 XOR2_X1 _5112_ (.A(_1361_),
    .B(_1371_),
    .Z(_1372_));
 XNOR2_X1 _5113_ (.A(_1359_),
    .B(_1372_),
    .ZN(_1373_));
 XOR2_X1 _5114_ (.A(_1357_),
    .B(_1373_),
    .Z(_1375_));
 XNOR2_X1 _5115_ (.A(_1356_),
    .B(_1375_),
    .ZN(_1376_));
 INV_X1 _5116_ (.A(_1312_),
    .ZN(_1377_));
 NAND2_X1 _5117_ (.A1(_1282_),
    .A2(_1377_),
    .ZN(_1378_));
 OR2_X1 _5118_ (.A1(_1284_),
    .A2(_1311_),
    .ZN(_1379_));
 AOI21_X1 _5119_ (.A(_1376_),
    .B1(_1378_),
    .B2(_1379_),
    .ZN(_1380_));
 AND3_X1 _5120_ (.A1(_1379_),
    .A2(_1378_),
    .A3(_1376_),
    .ZN(_1381_));
 NOR2_X1 _5121_ (.A1(_1380_),
    .A2(_1381_),
    .ZN(_1382_));
 XOR2_X1 _5122_ (.A(_1355_),
    .B(_1382_),
    .Z(_1383_));
 XNOR2_X1 _5123_ (.A(_0919_),
    .B(_1383_),
    .ZN(_1384_));
 XNOR2_X1 _5124_ (.A(_1354_),
    .B(_1384_),
    .ZN(_1386_));
 XNOR2_X1 _5125_ (.A(_1353_),
    .B(_1386_),
    .ZN(_1387_));
 OR2_X1 _5126_ (.A1(_1561_),
    .A2(_1323_),
    .ZN(_1388_));
 NAND2_X1 _5127_ (.A1(_1279_),
    .A2(_1322_),
    .ZN(_1389_));
 AOI21_X1 _5128_ (.A(_1387_),
    .B1(_1388_),
    .B2(_1389_),
    .ZN(_1390_));
 AND3_X1 _5129_ (.A1(_1389_),
    .A2(_1388_),
    .A3(_1387_),
    .ZN(_1391_));
 OR2_X1 _5130_ (.A1(_1390_),
    .A2(_1391_),
    .ZN(_1392_));
 OR2_X1 _5131_ (.A1(_0005_),
    .A2(_2731_),
    .ZN(_1393_));
 AOI21_X1 _5132_ (.A(_1392_),
    .B1(_1393_),
    .B2(_2586_),
    .ZN(_1394_));
 AND3_X1 _5133_ (.A1(_2586_),
    .A2(_1393_),
    .A3(_1392_),
    .ZN(_1395_));
 OR2_X1 _5134_ (.A1(_1394_),
    .A2(_1395_),
    .ZN(_1397_));
 XOR2_X1 _5135_ (.A(_1351_),
    .B(_1397_),
    .Z(_1398_));
 XNOR2_X1 _5136_ (.A(_1348_),
    .B(_1398_),
    .ZN(_1399_));
 NAND2_X1 _5137_ (.A1(_1347_),
    .A2(_1399_),
    .ZN(_1400_));
 XNOR2_X1 _5138_ (.A(_1347_),
    .B(_1399_),
    .ZN(_1401_));
 OAI21_X1 _5139_ (.A(_1328_),
    .B1(\coll_reg[10] ),
    .B2(\coll_reg[9] ),
    .ZN(_1402_));
 XOR2_X1 _5140_ (.A(_1402_),
    .B(_1344_),
    .Z(_1403_));
 NOR2_X1 _5141_ (.A1(\coll_reg[8] ),
    .A2(\coll_reg[10] ),
    .ZN(_1404_));
 NOR2_X1 _5142_ (.A1(_2659_),
    .A2(_1404_),
    .ZN(_1405_));
 XNOR2_X1 _5143_ (.A(\coll_reg[0] ),
    .B(_1331_),
    .ZN(_1406_));
 OR2_X1 _5144_ (.A1(_0919_),
    .A2(_1406_),
    .ZN(_1408_));
 XNOR2_X1 _5145_ (.A(\coll_reg[1] ),
    .B(_1333_),
    .ZN(_1409_));
 NOR2_X1 _5146_ (.A1(_1408_),
    .A2(_1409_),
    .ZN(_1410_));
 XOR2_X1 _5147_ (.A(_1408_),
    .B(_1409_),
    .Z(_1411_));
 AOI21_X1 _5148_ (.A(_1410_),
    .B1(_1411_),
    .B2(\coll_reg[5] ),
    .ZN(_1412_));
 XNOR2_X1 _5149_ (.A(\coll_reg[6] ),
    .B(_1339_),
    .ZN(_1413_));
 XOR2_X1 _5150_ (.A(_1412_),
    .B(_1413_),
    .Z(_1414_));
 NAND2_X1 _5151_ (.A1(_1405_),
    .A2(_1414_),
    .ZN(_1415_));
 OR2_X1 _5152_ (.A1(_1412_),
    .A2(_1413_),
    .ZN(_1416_));
 AOI21_X1 _5153_ (.A(_1403_),
    .B1(_1415_),
    .B2(_1416_),
    .ZN(_1417_));
 AND3_X1 _5154_ (.A1(_1346_),
    .A2(_1345_),
    .A3(_1327_),
    .ZN(_1419_));
 NOR2_X1 _5155_ (.A1(_1347_),
    .A2(_1419_),
    .ZN(_1420_));
 OR2_X1 _5156_ (.A1(_1417_),
    .A2(_1420_),
    .ZN(_1421_));
 AND2_X1 _5157_ (.A1(_1417_),
    .A2(_1420_),
    .ZN(_1422_));
 XNOR2_X1 _5158_ (.A(_1405_),
    .B(_1414_),
    .ZN(_1423_));
 XOR2_X1 _5159_ (.A(_1127_),
    .B(_1128_),
    .Z(_1424_));
 NAND2_X1 _5160_ (.A1(\coll_reg[3] ),
    .A2(_1424_),
    .ZN(_1425_));
 XNOR2_X1 _5161_ (.A(_0919_),
    .B(_1406_),
    .ZN(_1426_));
 NOR2_X1 _5162_ (.A1(_1425_),
    .A2(_1426_),
    .ZN(_1427_));
 XOR2_X1 _5163_ (.A(_1425_),
    .B(_1426_),
    .Z(_1428_));
 AOI21_X1 _5164_ (.A(_1427_),
    .B1(_1428_),
    .B2(\coll_reg[6] ),
    .ZN(_1430_));
 XNOR2_X1 _5165_ (.A(\coll_reg[5] ),
    .B(_1411_),
    .ZN(_1431_));
 XOR2_X1 _5166_ (.A(_1430_),
    .B(_1431_),
    .Z(_1432_));
 NAND2_X1 _5167_ (.A1(\coll_reg[7] ),
    .A2(_1432_),
    .ZN(_1433_));
 OR2_X1 _5168_ (.A1(_1430_),
    .A2(_1431_),
    .ZN(_1434_));
 AOI21_X1 _5169_ (.A(_1423_),
    .B1(_1433_),
    .B2(_1434_),
    .ZN(_1435_));
 AND3_X1 _5170_ (.A1(_1416_),
    .A2(_1415_),
    .A3(_1403_),
    .ZN(_1436_));
 NOR2_X1 _5171_ (.A1(_1417_),
    .A2(_1436_),
    .ZN(_1437_));
 NAND2_X1 _5172_ (.A1(_1435_),
    .A2(_1437_),
    .ZN(_1438_));
 NAND2_X1 _5173_ (.A1(_1434_),
    .A2(_1433_),
    .ZN(_1439_));
 XNOR2_X1 _5174_ (.A(_1439_),
    .B(_1423_),
    .ZN(_1441_));
 NOR3_X1 _5175_ (.A1(_0000_),
    .A2(_0007_),
    .A3(_2344_),
    .ZN(_1442_));
 XNOR2_X1 _5176_ (.A(\coll_reg[3] ),
    .B(_1424_),
    .ZN(_1443_));
 XNOR2_X1 _5177_ (.A(_1122_),
    .B(_1099_),
    .ZN(_1444_));
 XNOR2_X1 _5178_ (.A(_1125_),
    .B(_1444_),
    .ZN(_1445_));
 NAND2_X1 _5179_ (.A1(\coll_reg[1] ),
    .A2(_1445_),
    .ZN(_1446_));
 XOR2_X1 _5180_ (.A(_1098_),
    .B(_1126_),
    .Z(_1447_));
 XNOR2_X1 _5181_ (.A(_1446_),
    .B(_1447_),
    .ZN(_1448_));
 NAND3_X1 _5182_ (.A1(_2343_),
    .A2(_2344_),
    .A3(_1448_),
    .ZN(_1449_));
 NAND3_X1 _5183_ (.A1(\coll_reg[1] ),
    .A2(_1445_),
    .A3(_1447_),
    .ZN(_1450_));
 AOI21_X1 _5184_ (.A(_1443_),
    .B1(_1449_),
    .B2(_1450_),
    .ZN(_1452_));
 AND3_X1 _5185_ (.A1(_1450_),
    .A2(_1449_),
    .A3(_1443_),
    .ZN(_1453_));
 NOR2_X1 _5186_ (.A1(_1452_),
    .A2(_1453_),
    .ZN(_1454_));
 XOR2_X1 _5187_ (.A(_0007_),
    .B(_2344_),
    .Z(_1455_));
 AOI21_X1 _5188_ (.A(_1452_),
    .B1(_1454_),
    .B2(_1455_),
    .ZN(_1456_));
 XNOR2_X1 _5189_ (.A(\coll_reg[6] ),
    .B(_1428_),
    .ZN(_1457_));
 OR2_X1 _5190_ (.A1(_1456_),
    .A2(_1457_),
    .ZN(_1458_));
 XOR2_X1 _5191_ (.A(_1456_),
    .B(_1457_),
    .Z(_1459_));
 NOR2_X1 _5192_ (.A1(_0007_),
    .A2(_2344_),
    .ZN(_1460_));
 XNOR2_X1 _5193_ (.A(_0000_),
    .B(_1460_),
    .ZN(_1461_));
 NAND2_X1 _5194_ (.A1(_1459_),
    .A2(_1461_),
    .ZN(_1463_));
 NAND2_X1 _5195_ (.A1(_1458_),
    .A2(_1463_),
    .ZN(_1464_));
 XNOR2_X1 _5196_ (.A(\coll_reg[7] ),
    .B(_1432_),
    .ZN(_1465_));
 XNOR2_X1 _5197_ (.A(_1464_),
    .B(_1465_),
    .ZN(_1466_));
 AND2_X1 _5198_ (.A1(_1442_),
    .A2(_1466_),
    .ZN(_1467_));
 AOI21_X1 _5199_ (.A(_1465_),
    .B1(_1463_),
    .B2(_1458_),
    .ZN(_1468_));
 OAI21_X1 _5200_ (.A(_1441_),
    .B1(_1467_),
    .B2(_1468_),
    .ZN(_1469_));
 INV_X1 _5201_ (.A(_1469_),
    .ZN(_1470_));
 NOR2_X1 _5202_ (.A1(_1468_),
    .A2(_1467_),
    .ZN(_1471_));
 XNOR2_X1 _5203_ (.A(_1471_),
    .B(_1441_),
    .ZN(_1472_));
 XNOR2_X1 _5204_ (.A(_1454_),
    .B(_1455_),
    .ZN(_1474_));
 XNOR2_X1 _5205_ (.A(_2345_),
    .B(_1448_),
    .ZN(_1475_));
 XOR2_X1 _5206_ (.A(_1117_),
    .B(_1124_),
    .Z(_1476_));
 NAND2_X1 _5207_ (.A1(\coll_reg[0] ),
    .A2(_1476_),
    .ZN(_1477_));
 XNOR2_X1 _5208_ (.A(\coll_reg[1] ),
    .B(_1445_),
    .ZN(_1478_));
 XOR2_X1 _5209_ (.A(_1477_),
    .B(_1478_),
    .Z(_1479_));
 AND2_X1 _5210_ (.A1(\coll_reg[3] ),
    .A2(_1479_),
    .ZN(_1480_));
 NOR2_X1 _5211_ (.A1(_1477_),
    .A2(_1478_),
    .ZN(_1481_));
 OAI21_X1 _5212_ (.A(_1475_),
    .B1(_1480_),
    .B2(_1481_),
    .ZN(_1482_));
 OR3_X1 _5213_ (.A1(_1481_),
    .A2(_1480_),
    .A3(_1475_),
    .ZN(_1483_));
 AND2_X1 _5214_ (.A1(_1482_),
    .A2(_1483_),
    .ZN(_1485_));
 NAND2_X1 _5215_ (.A1(\coll_reg[7] ),
    .A2(_1485_),
    .ZN(_1486_));
 AOI21_X1 _5216_ (.A(_1474_),
    .B1(_1486_),
    .B2(_1482_),
    .ZN(_1487_));
 AND3_X1 _5217_ (.A1(_1482_),
    .A2(_1486_),
    .A3(_1474_),
    .ZN(_1488_));
 NOR2_X1 _5218_ (.A1(_1487_),
    .A2(_1488_),
    .ZN(_1489_));
 AOI21_X1 _5219_ (.A(_1487_),
    .B1(_1489_),
    .B2(\coll_reg[8] ),
    .ZN(_1490_));
 XNOR2_X1 _5220_ (.A(_1459_),
    .B(_1461_),
    .ZN(_1491_));
 NOR2_X1 _5221_ (.A1(_1490_),
    .A2(_1491_),
    .ZN(_1492_));
 XOR2_X1 _5222_ (.A(_1442_),
    .B(_1466_),
    .Z(_1493_));
 AND2_X1 _5223_ (.A1(_1492_),
    .A2(_1493_),
    .ZN(_1494_));
 XOR2_X1 _5224_ (.A(_1492_),
    .B(_1493_),
    .Z(_1496_));
 XNOR2_X1 _5225_ (.A(\coll_reg[7] ),
    .B(_1485_),
    .ZN(_1497_));
 XOR2_X1 _5226_ (.A(_1108_),
    .B(_1116_),
    .Z(_1498_));
 NAND2_X1 _5227_ (.A1(\coll_reg[1] ),
    .A2(_1498_),
    .ZN(_1499_));
 XNOR2_X1 _5228_ (.A(\coll_reg[0] ),
    .B(_1476_),
    .ZN(_1500_));
 NOR2_X1 _5229_ (.A1(_1499_),
    .A2(_1500_),
    .ZN(_1501_));
 XOR2_X1 _5230_ (.A(_1499_),
    .B(_1500_),
    .Z(_1502_));
 AOI21_X1 _5231_ (.A(_1501_),
    .B1(_1502_),
    .B2(\coll_reg[2] ),
    .ZN(_1503_));
 XNOR2_X1 _5232_ (.A(\coll_reg[3] ),
    .B(_1479_),
    .ZN(_1504_));
 XOR2_X1 _5233_ (.A(_1503_),
    .B(_1504_),
    .Z(_1505_));
 NAND2_X1 _5234_ (.A1(\coll_reg[6] ),
    .A2(_1505_),
    .ZN(_1507_));
 OR2_X1 _5235_ (.A1(_1503_),
    .A2(_1504_),
    .ZN(_1508_));
 AOI21_X1 _5236_ (.A(_1497_),
    .B1(_1507_),
    .B2(_1508_),
    .ZN(_1509_));
 XNOR2_X1 _5237_ (.A(_2585_),
    .B(_1489_),
    .ZN(_1510_));
 XOR2_X1 _5238_ (.A(_1490_),
    .B(_1491_),
    .Z(_1511_));
 NAND3_X1 _5239_ (.A1(_1509_),
    .A2(_1510_),
    .A3(_1511_),
    .ZN(_1512_));
 NAND2_X1 _5240_ (.A1(_1509_),
    .A2(_1510_),
    .ZN(_1513_));
 XNOR2_X1 _5241_ (.A(_1513_),
    .B(_1511_),
    .ZN(_1514_));
 XNOR2_X1 _5242_ (.A(\coll_reg[6] ),
    .B(_1505_),
    .ZN(_1515_));
 XOR2_X1 _5243_ (.A(_1103_),
    .B(_1107_),
    .Z(_1516_));
 XNOR2_X1 _5244_ (.A(\section_1.xn2[0] ),
    .B(_1516_),
    .ZN(_1518_));
 XNOR2_X1 _5245_ (.A(\coll_reg[1] ),
    .B(_1498_),
    .ZN(_1519_));
 NOR3_X1 _5246_ (.A1(_0749_),
    .A2(_1518_),
    .A3(_1519_),
    .ZN(_1520_));
 NOR2_X1 _5247_ (.A1(_0749_),
    .A2(_1518_),
    .ZN(_1521_));
 XNOR2_X1 _5248_ (.A(_1521_),
    .B(_1519_),
    .ZN(_1522_));
 AOI21_X1 _5249_ (.A(_1520_),
    .B1(_1522_),
    .B2(\coll_reg[4] ),
    .ZN(_1523_));
 XNOR2_X1 _5250_ (.A(\coll_reg[2] ),
    .B(_1502_),
    .ZN(_1524_));
 XOR2_X1 _5251_ (.A(_1523_),
    .B(_1524_),
    .Z(_1525_));
 NAND2_X1 _5252_ (.A1(\coll_reg[5] ),
    .A2(_1525_),
    .ZN(_1526_));
 OR2_X1 _5253_ (.A1(_1523_),
    .A2(_1524_),
    .ZN(_1527_));
 AOI21_X1 _5254_ (.A(_1515_),
    .B1(_1526_),
    .B2(_1527_),
    .ZN(_1529_));
 NAND2_X1 _5255_ (.A1(_1508_),
    .A2(_1507_),
    .ZN(_1530_));
 XNOR2_X1 _5256_ (.A(_1530_),
    .B(_1497_),
    .ZN(_1531_));
 AND2_X1 _5257_ (.A1(_1529_),
    .A2(_1531_),
    .ZN(_1532_));
 AND2_X1 _5258_ (.A1(_1510_),
    .A2(_1532_),
    .ZN(_1533_));
 XNOR2_X1 _5259_ (.A(_0749_),
    .B(_1518_),
    .ZN(_1534_));
 OR2_X1 _5260_ (.A1(_1286_),
    .A2(_1534_),
    .ZN(_1535_));
 XNOR2_X1 _5261_ (.A(\coll_reg[4] ),
    .B(_1522_),
    .ZN(_1536_));
 NOR2_X1 _5262_ (.A1(_1535_),
    .A2(_1536_),
    .ZN(_1537_));
 XNOR2_X1 _5263_ (.A(\coll_reg[5] ),
    .B(_1525_),
    .ZN(_1538_));
 INV_X1 _5264_ (.A(_1538_),
    .ZN(_1540_));
 NAND2_X1 _5265_ (.A1(_1527_),
    .A2(_1526_),
    .ZN(_1541_));
 XNOR2_X1 _5266_ (.A(_1541_),
    .B(_1515_),
    .ZN(_1542_));
 NAND3_X1 _5267_ (.A1(_1537_),
    .A2(_1540_),
    .A3(_1542_),
    .ZN(_1543_));
 XNOR2_X1 _5268_ (.A(_1529_),
    .B(_1531_),
    .ZN(_1544_));
 XOR2_X1 _5269_ (.A(_1543_),
    .B(_1544_),
    .Z(_1545_));
 XNOR2_X1 _5270_ (.A(_1286_),
    .B(_1534_),
    .ZN(_1546_));
 NAND2_X1 _5271_ (.A1(\coll_reg[1] ),
    .A2(\section_1.t1[1] ),
    .ZN(_1547_));
 XNOR2_X1 _5272_ (.A(\section_1.xn2[0] ),
    .B(_1102_),
    .ZN(_1548_));
 XOR2_X1 _5273_ (.A(_1547_),
    .B(_1548_),
    .Z(_1549_));
 NAND2_X1 _5274_ (.A1(\coll_reg[2] ),
    .A2(_1549_),
    .ZN(_1551_));
 OR2_X1 _5275_ (.A1(_1547_),
    .A2(_1548_),
    .ZN(_1552_));
 AOI21_X1 _5276_ (.A(_1546_),
    .B1(_1551_),
    .B2(_1552_),
    .ZN(_1553_));
 XOR2_X1 _5277_ (.A(_1535_),
    .B(_1536_),
    .Z(_1554_));
 AND3_X1 _5278_ (.A1(_1540_),
    .A2(_1553_),
    .A3(_1554_),
    .ZN(_1555_));
 NAND2_X1 _5279_ (.A1(_1537_),
    .A2(_1540_),
    .ZN(_1556_));
 XNOR2_X1 _5280_ (.A(_1556_),
    .B(_1542_),
    .ZN(_1557_));
 NAND2_X1 _5281_ (.A1(_1555_),
    .A2(_1557_),
    .ZN(_1558_));
 XOR2_X1 _5282_ (.A(\coll_reg[1] ),
    .B(\section_1.t1[1] ),
    .Z(_1559_));
 NAND3_X1 _5283_ (.A1(\coll_reg[0] ),
    .A2(\section_1.t1[0] ),
    .A3(_1559_),
    .ZN(_1560_));
 XNOR2_X1 _5284_ (.A(\coll_reg[2] ),
    .B(_1549_),
    .ZN(_1562_));
 NOR2_X1 _5285_ (.A1(_1560_),
    .A2(_1562_),
    .ZN(_1563_));
 AND3_X1 _5286_ (.A1(_1552_),
    .A2(_1551_),
    .A3(_1546_),
    .ZN(_1564_));
 NOR2_X1 _5287_ (.A1(_1553_),
    .A2(_1564_),
    .ZN(_1565_));
 NAND2_X1 _5288_ (.A1(_1563_),
    .A2(_1565_),
    .ZN(_1566_));
 XNOR2_X1 _5289_ (.A(_1553_),
    .B(_1554_),
    .ZN(_1567_));
 OR2_X1 _5290_ (.A1(_1566_),
    .A2(_1567_),
    .ZN(_1568_));
 AOI21_X1 _5291_ (.A(_1537_),
    .B1(_1553_),
    .B2(_1554_),
    .ZN(_1569_));
 XNOR2_X1 _5292_ (.A(_1538_),
    .B(_1569_),
    .ZN(_1570_));
 OR2_X1 _5293_ (.A1(_1568_),
    .A2(_1570_),
    .ZN(_1571_));
 XNOR2_X1 _5294_ (.A(_1555_),
    .B(_1557_),
    .ZN(_1573_));
 OAI21_X1 _5295_ (.A(_1558_),
    .B1(_1571_),
    .B2(_1573_),
    .ZN(_1574_));
 NAND2_X1 _5296_ (.A1(_1545_),
    .A2(_1574_),
    .ZN(_1575_));
 OAI21_X1 _5297_ (.A(_1575_),
    .B1(_1544_),
    .B2(_1543_),
    .ZN(_1576_));
 NOR2_X1 _5298_ (.A1(_1509_),
    .A2(_1532_),
    .ZN(_1577_));
 XNOR2_X1 _5299_ (.A(_1510_),
    .B(_1577_),
    .ZN(_1578_));
 AND2_X1 _5300_ (.A1(_1576_),
    .A2(_1578_),
    .ZN(_1579_));
 OAI21_X1 _5301_ (.A(_1514_),
    .B1(_1533_),
    .B2(_1579_),
    .ZN(_1580_));
 NAND2_X1 _5302_ (.A1(_1512_),
    .A2(_1580_),
    .ZN(_1581_));
 AOI21_X1 _5303_ (.A(_1494_),
    .B1(_1496_),
    .B2(_1581_),
    .ZN(_1582_));
 INV_X1 _5304_ (.A(_1582_),
    .ZN(_1584_));
 AOI21_X1 _5305_ (.A(_1470_),
    .B1(_1472_),
    .B2(_1584_),
    .ZN(_1585_));
 XNOR2_X1 _5306_ (.A(_1435_),
    .B(_1437_),
    .ZN(_1586_));
 OAI21_X1 _5307_ (.A(_1438_),
    .B1(_1585_),
    .B2(_1586_),
    .ZN(_1587_));
 OAI21_X1 _5308_ (.A(_1421_),
    .B1(_1422_),
    .B2(_1587_),
    .ZN(_1588_));
 OAI21_X1 _5309_ (.A(_1400_),
    .B1(_1401_),
    .B2(_1588_),
    .ZN(_1589_));
 AOI21_X1 _5310_ (.A(_1397_),
    .B1(_1350_),
    .B2(_1349_),
    .ZN(_1590_));
 NOR4_X1 _5311_ (.A1(\coll_reg[9] ),
    .A2(_0005_),
    .A3(_2732_),
    .A4(_1398_),
    .ZN(_1591_));
 OR2_X1 _5312_ (.A1(_1590_),
    .A2(_1591_),
    .ZN(_1592_));
 NAND4_X1 _5313_ (.A1(\coll_reg[9] ),
    .A2(\coll_reg[5] ),
    .A3(\coll_reg[10] ),
    .A4(_1924_),
    .ZN(_1593_));
 OAI21_X1 _5314_ (.A(_2731_),
    .B1(_2282_),
    .B2(_2283_),
    .ZN(_1595_));
 NAND2_X1 _5315_ (.A1(_1593_),
    .A2(_1595_),
    .ZN(_1596_));
 NAND2_X1 _5316_ (.A1(_1354_),
    .A2(_1384_),
    .ZN(_1597_));
 OAI21_X1 _5317_ (.A(_1597_),
    .B1(_1386_),
    .B2(_1353_),
    .ZN(_1598_));
 AND2_X1 _5318_ (.A1(\coll_reg[4] ),
    .A2(_1383_),
    .ZN(_1599_));
 NAND2_X1 _5319_ (.A1(\section_1.xn2[9] ),
    .A2(_1296_),
    .ZN(_1600_));
 NAND2_X1 _5320_ (.A1(_0933_),
    .A2(\section_1.xn2[10] ),
    .ZN(_1601_));
 NAND2_X1 _5321_ (.A1(_1362_),
    .A2(_1370_),
    .ZN(_1602_));
 OAI21_X1 _5322_ (.A(_1602_),
    .B1(_1369_),
    .B2(_0010_),
    .ZN(_1603_));
 NAND3_X1 _5323_ (.A1(_0920_),
    .A2(_0921_),
    .A3(_0922_),
    .ZN(_1604_));
 OAI21_X1 _5324_ (.A(\section_1.xn1[10] ),
    .B1(_1604_),
    .B2(\section_1.xn1[6] ),
    .ZN(_1606_));
 NAND2_X1 _5325_ (.A1(_1368_),
    .A2(_1606_),
    .ZN(_1607_));
 XNOR2_X1 _5326_ (.A(_1364_),
    .B(_1607_),
    .ZN(_1608_));
 XNOR2_X1 _5327_ (.A(_1362_),
    .B(_1608_),
    .ZN(_1609_));
 XOR2_X1 _5328_ (.A(_1603_),
    .B(_1609_),
    .Z(_1610_));
 XNOR2_X1 _5329_ (.A(_1601_),
    .B(_1610_),
    .ZN(_1611_));
 AND2_X1 _5330_ (.A1(_1359_),
    .A2(_1372_),
    .ZN(_1612_));
 NOR2_X1 _5331_ (.A1(_1361_),
    .A2(_1371_),
    .ZN(_1613_));
 OAI21_X1 _5332_ (.A(_1611_),
    .B1(_1612_),
    .B2(_1613_),
    .ZN(_1614_));
 OR3_X1 _5333_ (.A1(_1613_),
    .A2(_1612_),
    .A3(_1611_),
    .ZN(_1615_));
 AND2_X1 _5334_ (.A1(_1614_),
    .A2(_1615_),
    .ZN(_1617_));
 XNOR2_X1 _5335_ (.A(_1600_),
    .B(_1617_),
    .ZN(_1618_));
 AND2_X1 _5336_ (.A1(_1356_),
    .A2(_1375_),
    .ZN(_1619_));
 NOR2_X1 _5337_ (.A1(_1357_),
    .A2(_1373_),
    .ZN(_1620_));
 OAI21_X1 _5338_ (.A(_1618_),
    .B1(_1619_),
    .B2(_1620_),
    .ZN(_1621_));
 OR3_X1 _5339_ (.A1(_1620_),
    .A2(_1619_),
    .A3(_1618_),
    .ZN(_1622_));
 AND2_X1 _5340_ (.A1(_1621_),
    .A2(_1622_),
    .ZN(_1623_));
 AND2_X1 _5341_ (.A1(_1355_),
    .A2(_1382_),
    .ZN(_1624_));
 NOR2_X1 _5342_ (.A1(_1380_),
    .A2(_1624_),
    .ZN(_1625_));
 XNOR2_X1 _5343_ (.A(_1623_),
    .B(_1625_),
    .ZN(_1626_));
 XOR2_X1 _5344_ (.A(_1599_),
    .B(_1626_),
    .Z(_1628_));
 XOR2_X1 _5345_ (.A(_2285_),
    .B(_1628_),
    .Z(_1629_));
 XNOR2_X1 _5346_ (.A(_1598_),
    .B(_1629_),
    .ZN(_1630_));
 XOR2_X1 _5347_ (.A(_1596_),
    .B(_1630_),
    .Z(_1631_));
 OAI21_X1 _5348_ (.A(_1631_),
    .B1(_1394_),
    .B2(_1390_),
    .ZN(_1632_));
 OR3_X1 _5349_ (.A1(_1390_),
    .A2(_1394_),
    .A3(_1631_),
    .ZN(_1633_));
 AND2_X1 _5350_ (.A1(_1632_),
    .A2(_1633_),
    .ZN(_1634_));
 XOR2_X1 _5351_ (.A(_1592_),
    .B(_1634_),
    .Z(_1635_));
 XNOR2_X1 _5352_ (.A(_1589_),
    .B(_1635_),
    .ZN(_1636_));
 XNOR2_X1 _5353_ (.A(_2717_),
    .B(_1636_),
    .ZN(_1637_));
 XOR2_X1 _5354_ (.A(\section_1.yn2[9] ),
    .B(\section_1.yn2[10] ),
    .Z(_1639_));
 XOR2_X1 _5355_ (.A(_1401_),
    .B(_1588_),
    .Z(_1640_));
 XNOR2_X1 _5356_ (.A(_0004_),
    .B(_1640_),
    .ZN(_1641_));
 NAND2_X1 _5357_ (.A1(_1639_),
    .A2(_1641_),
    .ZN(_1642_));
 NAND2_X1 _5358_ (.A1(_0144_),
    .A2(_1640_),
    .ZN(_1643_));
 AOI21_X1 _5359_ (.A(_1637_),
    .B1(_1642_),
    .B2(_1643_),
    .ZN(_1644_));
 XNOR2_X1 _5360_ (.A(_0938_),
    .B(_0940_),
    .ZN(_1645_));
 AND3_X1 _5361_ (.A1(_1643_),
    .A2(_1642_),
    .A3(_1637_),
    .ZN(_1646_));
 OR2_X1 _5362_ (.A1(_1644_),
    .A2(_1646_),
    .ZN(_1647_));
 NOR2_X1 _5363_ (.A1(_1645_),
    .A2(_1647_),
    .ZN(_1648_));
 NOR2_X1 _5364_ (.A1(_1644_),
    .A2(_1648_),
    .ZN(_1650_));
 INV_X1 _5365_ (.A(_1650_),
    .ZN(_1651_));
 NAND2_X1 _5366_ (.A1(\section_1.yn2[9] ),
    .A2(\section_1.yn2[7] ),
    .ZN(_1652_));
 XNOR2_X1 _5367_ (.A(_2504_),
    .B(_1652_),
    .ZN(_1653_));
 XNOR2_X1 _5368_ (.A(\section_1.yn2[10] ),
    .B(_0004_),
    .ZN(_1654_));
 XNOR2_X1 _5369_ (.A(_1636_),
    .B(_1654_),
    .ZN(_1655_));
 NAND2_X1 _5370_ (.A1(_0144_),
    .A2(_1655_),
    .ZN(_1656_));
 NAND2_X1 _5371_ (.A1(_1592_),
    .A2(_1634_),
    .ZN(_1657_));
 NAND2_X1 _5372_ (.A1(_1589_),
    .A2(_1635_),
    .ZN(_1658_));
 NAND2_X1 _5373_ (.A1(_1657_),
    .A2(_1658_),
    .ZN(_1659_));
 NAND2_X1 _5374_ (.A1(_1598_),
    .A2(_1629_),
    .ZN(_1661_));
 OAI21_X1 _5375_ (.A(_1661_),
    .B1(_1630_),
    .B2(_1596_),
    .ZN(_1662_));
 NAND2_X1 _5376_ (.A1(_1624_),
    .A2(_1623_),
    .ZN(_1663_));
 NAND2_X1 _5377_ (.A1(_1380_),
    .A2(_1622_),
    .ZN(_1664_));
 NAND3_X1 _5378_ (.A1(_1621_),
    .A2(_1663_),
    .A3(_1664_),
    .ZN(_1665_));
 NAND2_X1 _5379_ (.A1(\in_reg1[10] ),
    .A2(\section_1.xn2[10] ),
    .ZN(_1666_));
 NAND2_X1 _5380_ (.A1(_1603_),
    .A2(_1609_),
    .ZN(_1667_));
 INV_X1 _5381_ (.A(_1610_),
    .ZN(_1668_));
 OAI21_X1 _5382_ (.A(_1667_),
    .B1(_1668_),
    .B2(_1601_),
    .ZN(_1669_));
 XNOR2_X1 _5383_ (.A(\section_1.xn1[10] ),
    .B(_0010_),
    .ZN(_1670_));
 XNOR2_X1 _5384_ (.A(_1362_),
    .B(_1670_),
    .ZN(_1672_));
 INV_X1 _5385_ (.A(_1608_),
    .ZN(_1673_));
 NAND2_X1 _5386_ (.A1(_1362_),
    .A2(_1673_),
    .ZN(_1674_));
 NAND2_X1 _5387_ (.A1(_1364_),
    .A2(_1607_),
    .ZN(_1675_));
 AOI21_X1 _5388_ (.A(_1672_),
    .B1(_1674_),
    .B2(_1675_),
    .ZN(_1676_));
 AND3_X1 _5389_ (.A1(_1675_),
    .A2(_1674_),
    .A3(_1672_),
    .ZN(_1677_));
 OR2_X1 _5390_ (.A1(_1676_),
    .A2(_1677_),
    .ZN(_1678_));
 XOR2_X1 _5391_ (.A(_1601_),
    .B(_1678_),
    .Z(_1679_));
 XNOR2_X1 _5392_ (.A(_1669_),
    .B(_1679_),
    .ZN(_1680_));
 XNOR2_X1 _5393_ (.A(_1666_),
    .B(_1680_),
    .ZN(_1681_));
 NAND3_X1 _5394_ (.A1(\section_1.xn2[9] ),
    .A2(_1296_),
    .A3(_1617_),
    .ZN(_1683_));
 AOI21_X1 _5395_ (.A(_1681_),
    .B1(_1683_),
    .B2(_1614_),
    .ZN(_1684_));
 AND3_X1 _5396_ (.A1(_1614_),
    .A2(_1683_),
    .A3(_1681_),
    .ZN(_1685_));
 NOR2_X1 _5397_ (.A1(_1684_),
    .A2(_1685_),
    .ZN(_1686_));
 XNOR2_X1 _5398_ (.A(_1665_),
    .B(_1686_),
    .ZN(_1687_));
 NAND2_X1 _5399_ (.A1(\coll_reg[6] ),
    .A2(\coll_reg[5] ),
    .ZN(_1688_));
 XNOR2_X1 _5400_ (.A(_1688_),
    .B(_2340_),
    .ZN(_1689_));
 XOR2_X1 _5401_ (.A(_1687_),
    .B(_1689_),
    .Z(_1690_));
 NAND2_X1 _5402_ (.A1(_2285_),
    .A2(_1628_),
    .ZN(_1691_));
 NAND2_X1 _5403_ (.A1(_1599_),
    .A2(_1626_),
    .ZN(_1692_));
 AOI21_X1 _5404_ (.A(_1690_),
    .B1(_1691_),
    .B2(_1692_),
    .ZN(_1694_));
 AND3_X1 _5405_ (.A1(_1692_),
    .A2(_1691_),
    .A3(_1690_),
    .ZN(_1695_));
 OR2_X1 _5406_ (.A1(_1694_),
    .A2(_1695_),
    .ZN(_1696_));
 XNOR2_X1 _5407_ (.A(_0330_),
    .B(_1696_),
    .ZN(_1697_));
 XOR2_X1 _5408_ (.A(_1662_),
    .B(_1697_),
    .Z(_1698_));
 XNOR2_X1 _5409_ (.A(_1593_),
    .B(_1698_),
    .ZN(_1699_));
 XOR2_X1 _5410_ (.A(_1632_),
    .B(_1699_),
    .Z(_1700_));
 XOR2_X1 _5411_ (.A(_1659_),
    .B(_1700_),
    .Z(_1701_));
 XNOR2_X1 _5412_ (.A(\section_1.yn2[10] ),
    .B(_1701_),
    .ZN(_1702_));
 XOR2_X1 _5413_ (.A(_1656_),
    .B(_1702_),
    .Z(_1703_));
 XNOR2_X1 _5414_ (.A(_1653_),
    .B(_1703_),
    .ZN(_1705_));
 XOR2_X1 _5415_ (.A(_0003_),
    .B(_0941_),
    .Z(_1706_));
 XNOR2_X1 _5416_ (.A(_1650_),
    .B(_1705_),
    .ZN(_1707_));
 AOI22_X1 _5417_ (.A1(_1651_),
    .A2(_1705_),
    .B1(_1706_),
    .B2(_1707_),
    .ZN(_1708_));
 MUX2_X1 _5418_ (.A(_0004_),
    .B(_1652_),
    .S(\section_1.yn2[8] ),
    .Z(_1709_));
 XOR2_X1 _5419_ (.A(_0001_),
    .B(_1709_),
    .Z(_1710_));
 NOR2_X1 _5420_ (.A1(_1656_),
    .A2(_1702_),
    .ZN(_1711_));
 INV_X1 _5421_ (.A(_1653_),
    .ZN(_1712_));
 AOI21_X1 _5422_ (.A(_1711_),
    .B1(_1703_),
    .B2(_1712_),
    .ZN(_1713_));
 NAND2_X1 _5423_ (.A1(\section_1.yn2[8] ),
    .A2(\section_1.yn2[10] ),
    .ZN(_1714_));
 XNOR2_X1 _5424_ (.A(_2572_),
    .B(_1714_),
    .ZN(_1716_));
 XNOR2_X1 _5425_ (.A(_1654_),
    .B(_1701_),
    .ZN(_1717_));
 NOR2_X1 _5426_ (.A1(_0004_),
    .A2(_1717_),
    .ZN(_1718_));
 NOR2_X1 _5427_ (.A1(_1632_),
    .A2(_1699_),
    .ZN(_1719_));
 AOI21_X1 _5428_ (.A(_1719_),
    .B1(_1700_),
    .B2(_1659_),
    .ZN(_1720_));
 INV_X1 _5429_ (.A(_1697_),
    .ZN(_1721_));
 NAND2_X1 _5430_ (.A1(_1662_),
    .A2(_1721_),
    .ZN(_1722_));
 OAI21_X1 _5431_ (.A(_1722_),
    .B1(_1698_),
    .B2(_1593_),
    .ZN(_1723_));
 INV_X1 _5432_ (.A(_1696_),
    .ZN(_1724_));
 AOI21_X1 _5433_ (.A(_1694_),
    .B1(_1724_),
    .B2(\coll_reg[10] ),
    .ZN(_1725_));
 NOR2_X1 _5434_ (.A1(\coll_reg[7] ),
    .A2(_1688_),
    .ZN(_1727_));
 XOR2_X1 _5435_ (.A(_1405_),
    .B(_1727_),
    .Z(_1728_));
 INV_X1 _5436_ (.A(_1687_),
    .ZN(_1729_));
 NAND2_X1 _5437_ (.A1(_1729_),
    .A2(_1689_),
    .ZN(_1730_));
 NOR2_X1 _5438_ (.A1(_0918_),
    .A2(\coll_reg[6] ),
    .ZN(_1731_));
 AOI21_X1 _5439_ (.A(_1684_),
    .B1(_1686_),
    .B2(_1665_),
    .ZN(_1732_));
 NAND2_X1 _5440_ (.A1(_1669_),
    .A2(_1679_),
    .ZN(_1733_));
 OAI21_X1 _5441_ (.A(_1733_),
    .B1(_1680_),
    .B2(_1666_),
    .ZN(_1734_));
 NOR3_X1 _5442_ (.A1(\section_1.xn1[10] ),
    .A2(_1364_),
    .A3(_1362_),
    .ZN(_1735_));
 AOI21_X1 _5443_ (.A(_1601_),
    .B1(_1364_),
    .B2(\section_1.xn1[10] ),
    .ZN(_1736_));
 NAND2_X1 _5444_ (.A1(\in_reg1[10] ),
    .A2(_1285_),
    .ZN(_1738_));
 NOR3_X1 _5445_ (.A1(_0927_),
    .A2(_0010_),
    .A3(_1738_),
    .ZN(_1739_));
 NOR3_X1 _5446_ (.A1(_1735_),
    .A2(_1736_),
    .A3(_1739_),
    .ZN(_1740_));
 NOR2_X1 _5447_ (.A1(_1601_),
    .A2(_1678_),
    .ZN(_1741_));
 OAI21_X1 _5448_ (.A(_1740_),
    .B1(_1741_),
    .B2(_1676_),
    .ZN(_1742_));
 OR3_X1 _5449_ (.A1(_1676_),
    .A2(_1741_),
    .A3(_1740_),
    .ZN(_1743_));
 AND2_X1 _5450_ (.A1(_1742_),
    .A2(_1743_),
    .ZN(_1744_));
 XNOR2_X1 _5451_ (.A(_1666_),
    .B(_1744_),
    .ZN(_1745_));
 NAND2_X1 _5452_ (.A1(_1734_),
    .A2(_1745_),
    .ZN(_1746_));
 OR2_X1 _5453_ (.A1(_1734_),
    .A2(_1745_),
    .ZN(_1747_));
 AND3_X1 _5454_ (.A1(_1732_),
    .A2(_1746_),
    .A3(_1747_),
    .ZN(_1749_));
 XNOR2_X1 _5455_ (.A(_1731_),
    .B(_1749_),
    .ZN(_1750_));
 XOR2_X1 _5456_ (.A(_1730_),
    .B(_1750_),
    .Z(_1751_));
 XNOR2_X1 _5457_ (.A(_1728_),
    .B(_1751_),
    .ZN(_1752_));
 XOR2_X1 _5458_ (.A(_1725_),
    .B(_1752_),
    .Z(_1753_));
 XNOR2_X1 _5459_ (.A(_1723_),
    .B(_1753_),
    .ZN(_1754_));
 XNOR2_X1 _5460_ (.A(_1720_),
    .B(_1754_),
    .ZN(_1755_));
 XNOR2_X1 _5461_ (.A(\section_1.yn2[10] ),
    .B(_1755_),
    .ZN(_1756_));
 XNOR2_X1 _5462_ (.A(_1718_),
    .B(_1756_),
    .ZN(_1757_));
 XNOR2_X1 _5463_ (.A(_1716_),
    .B(_1757_),
    .ZN(_1758_));
 XNOR2_X1 _5464_ (.A(_1713_),
    .B(_1758_),
    .ZN(_1760_));
 XNOR2_X1 _5465_ (.A(_1710_),
    .B(_1760_),
    .ZN(_1761_));
 XOR2_X1 _5466_ (.A(_1708_),
    .B(_1761_),
    .Z(_1762_));
 NAND3_X1 _5467_ (.A1(_0003_),
    .A2(_0941_),
    .A3(_1762_),
    .ZN(_1763_));
 OAI21_X1 _5468_ (.A(_1763_),
    .B1(_1761_),
    .B2(_1708_),
    .ZN(_1764_));
 INV_X1 _5469_ (.A(_1709_),
    .ZN(_1765_));
 NAND2_X1 _5470_ (.A1(_0001_),
    .A2(_1765_),
    .ZN(_1766_));
 OAI22_X1 _5471_ (.A1(\section_1.yn2[9] ),
    .A2(_0004_),
    .B1(_0937_),
    .B2(_2504_),
    .ZN(_1767_));
 XOR2_X1 _5472_ (.A(_0008_),
    .B(_1767_),
    .Z(_1768_));
 NAND2_X1 _5473_ (.A1(_1718_),
    .A2(_1756_),
    .ZN(_1769_));
 OAI21_X1 _5474_ (.A(_1769_),
    .B1(_1757_),
    .B2(_1716_),
    .ZN(_1771_));
 NOR2_X1 _5475_ (.A1(\section_1.yn2[9] ),
    .A2(_2717_),
    .ZN(_1772_));
 XNOR2_X1 _5476_ (.A(_1654_),
    .B(_1755_),
    .ZN(_1773_));
 AND2_X1 _5477_ (.A1(_0144_),
    .A2(_1773_),
    .ZN(_1774_));
 AND2_X1 _5478_ (.A1(_1723_),
    .A2(_1753_),
    .ZN(_1775_));
 NOR2_X1 _5479_ (.A1(_1720_),
    .A2(_1754_),
    .ZN(_1776_));
 NOR2_X1 _5480_ (.A1(_1725_),
    .A2(_1752_),
    .ZN(_1777_));
 AND2_X1 _5481_ (.A1(_1405_),
    .A2(_1727_),
    .ZN(_1778_));
 NOR2_X1 _5482_ (.A1(_1730_),
    .A2(_1750_),
    .ZN(_1779_));
 AOI21_X1 _5483_ (.A(_1779_),
    .B1(_1751_),
    .B2(_1728_),
    .ZN(_1780_));
 AND2_X1 _5484_ (.A1(_2585_),
    .A2(_2586_),
    .ZN(_1782_));
 NOR2_X1 _5485_ (.A1(_2588_),
    .A2(_1782_),
    .ZN(_1783_));
 XNOR2_X1 _5486_ (.A(_2452_),
    .B(_1783_),
    .ZN(_1784_));
 INV_X1 _5487_ (.A(_1784_),
    .ZN(_1785_));
 AND2_X1 _5488_ (.A1(_1731_),
    .A2(_1749_),
    .ZN(_1786_));
 NAND2_X1 _5489_ (.A1(_1732_),
    .A2(_1746_),
    .ZN(_1787_));
 INV_X1 _5490_ (.A(_1744_),
    .ZN(_1788_));
 OAI21_X1 _5491_ (.A(_1742_),
    .B1(_1788_),
    .B2(_1666_),
    .ZN(_1789_));
 NAND3_X1 _5492_ (.A1(\section_1.xn1[10] ),
    .A2(_0010_),
    .A3(_1738_),
    .ZN(_1790_));
 NAND2_X1 _5493_ (.A1(_1601_),
    .A2(_1790_),
    .ZN(_1791_));
 OAI21_X1 _5494_ (.A(_1791_),
    .B1(_0010_),
    .B2(\section_1.xn1[10] ),
    .ZN(_1793_));
 OAI21_X1 _5495_ (.A(_1793_),
    .B1(_1738_),
    .B2(_0010_),
    .ZN(_1794_));
 XNOR2_X1 _5496_ (.A(_1789_),
    .B(_1794_),
    .ZN(_1795_));
 XNOR2_X1 _5497_ (.A(_1787_),
    .B(_1795_),
    .ZN(_1796_));
 XNOR2_X1 _5498_ (.A(_1786_),
    .B(_1796_),
    .ZN(_1797_));
 XNOR2_X1 _5499_ (.A(_1785_),
    .B(_1797_),
    .ZN(_1798_));
 XOR2_X1 _5500_ (.A(_1780_),
    .B(_1798_),
    .Z(_1799_));
 XOR2_X1 _5501_ (.A(_1778_),
    .B(_1799_),
    .Z(_1800_));
 XOR2_X1 _5502_ (.A(_1777_),
    .B(_1800_),
    .Z(_1801_));
 OR3_X1 _5503_ (.A1(_1775_),
    .A2(_1776_),
    .A3(_1801_),
    .ZN(_1802_));
 OAI21_X1 _5504_ (.A(_1801_),
    .B1(_1776_),
    .B2(_1775_),
    .ZN(_1804_));
 NAND2_X1 _5505_ (.A1(_1802_),
    .A2(_1804_),
    .ZN(_1805_));
 XNOR2_X1 _5506_ (.A(\section_1.yn2[10] ),
    .B(_1805_),
    .ZN(_1806_));
 XNOR2_X1 _5507_ (.A(_1774_),
    .B(_1806_),
    .ZN(_1807_));
 XNOR2_X1 _5508_ (.A(_1772_),
    .B(_1807_),
    .ZN(_1808_));
 XOR2_X1 _5509_ (.A(_1771_),
    .B(_1808_),
    .Z(_1809_));
 XOR2_X1 _5510_ (.A(_1768_),
    .B(_1809_),
    .Z(_1810_));
 NOR2_X1 _5511_ (.A1(_1710_),
    .A2(_1760_),
    .ZN(_1811_));
 NOR2_X1 _5512_ (.A1(_1713_),
    .A2(_1758_),
    .ZN(_1812_));
 OAI21_X1 _5513_ (.A(_1810_),
    .B1(_1811_),
    .B2(_1812_),
    .ZN(_1813_));
 OR3_X1 _5514_ (.A1(_1812_),
    .A2(_1811_),
    .A3(_1810_),
    .ZN(_1815_));
 NAND2_X1 _5515_ (.A1(_1813_),
    .A2(_1815_),
    .ZN(_1816_));
 XOR2_X1 _5516_ (.A(_1766_),
    .B(_1816_),
    .Z(_1817_));
 NAND2_X1 _5517_ (.A1(_1764_),
    .A2(_1817_),
    .ZN(_1818_));
 NOR2_X1 _5518_ (.A1(_1764_),
    .A2(_1817_),
    .ZN(_1819_));
 XOR2_X1 _5519_ (.A(_1417_),
    .B(_1420_),
    .Z(_1820_));
 XNOR2_X1 _5520_ (.A(_1587_),
    .B(_1820_),
    .ZN(_1821_));
 OR2_X1 _5521_ (.A1(_0004_),
    .A2(_1821_),
    .ZN(_1822_));
 XNOR2_X1 _5522_ (.A(\section_1.yn2[8] ),
    .B(\section_1.yn2[10] ),
    .ZN(_1823_));
 XNOR2_X1 _5523_ (.A(_0004_),
    .B(_1821_),
    .ZN(_1824_));
 OAI21_X1 _5524_ (.A(_1822_),
    .B1(_1823_),
    .B2(_1824_),
    .ZN(_1826_));
 XOR2_X1 _5525_ (.A(_1639_),
    .B(_1641_),
    .Z(_1827_));
 NAND2_X1 _5526_ (.A1(_1826_),
    .A2(_1827_),
    .ZN(_1828_));
 NAND2_X1 _5527_ (.A1(\section_1.yn2[7] ),
    .A2(\section_1.yn2[5] ),
    .ZN(_1829_));
 XOR2_X1 _5528_ (.A(\section_1.yn2[8] ),
    .B(\section_1.yn2[6] ),
    .Z(_1830_));
 XNOR2_X1 _5529_ (.A(_1714_),
    .B(_1830_),
    .ZN(_1831_));
 XNOR2_X1 _5530_ (.A(_1829_),
    .B(_1831_),
    .ZN(_1832_));
 INV_X1 _5531_ (.A(_1832_),
    .ZN(_1833_));
 XNOR2_X1 _5532_ (.A(_1826_),
    .B(_1827_),
    .ZN(_1834_));
 OAI21_X1 _5533_ (.A(_1828_),
    .B1(_1833_),
    .B2(_1834_),
    .ZN(_1835_));
 INV_X1 _5534_ (.A(_1835_),
    .ZN(_1837_));
 XNOR2_X1 _5535_ (.A(_1645_),
    .B(_1647_),
    .ZN(_1838_));
 NOR2_X1 _5536_ (.A1(_1837_),
    .A2(_1838_),
    .ZN(_1839_));
 NAND3_X1 _5537_ (.A1(\section_1.yn2[7] ),
    .A2(\section_1.yn2[5] ),
    .A3(_1831_),
    .ZN(_1840_));
 OAI21_X1 _5538_ (.A(_1840_),
    .B1(_1714_),
    .B2(\section_1.yn2[6] ),
    .ZN(_1841_));
 XOR2_X1 _5539_ (.A(_0009_),
    .B(_1841_),
    .Z(_1842_));
 XNOR2_X1 _5540_ (.A(_1835_),
    .B(_1838_),
    .ZN(_1843_));
 AOI21_X1 _5541_ (.A(_1839_),
    .B1(_1842_),
    .B2(_1843_),
    .ZN(_1844_));
 XNOR2_X1 _5542_ (.A(_1706_),
    .B(_1707_),
    .ZN(_1845_));
 OR2_X1 _5543_ (.A1(_1844_),
    .A2(_1845_),
    .ZN(_1846_));
 XNOR2_X1 _5544_ (.A(_1844_),
    .B(_1845_),
    .ZN(_1848_));
 NAND2_X1 _5545_ (.A1(_0009_),
    .A2(_1841_),
    .ZN(_1849_));
 OAI21_X1 _5546_ (.A(_1846_),
    .B1(_1848_),
    .B2(_1849_),
    .ZN(_1850_));
 NAND2_X1 _5547_ (.A1(_0003_),
    .A2(_0941_),
    .ZN(_1851_));
 XNOR2_X1 _5548_ (.A(_1851_),
    .B(_1762_),
    .ZN(_1852_));
 NAND2_X1 _5549_ (.A1(_1850_),
    .A2(_1852_),
    .ZN(_1853_));
 XOR2_X1 _5550_ (.A(_1850_),
    .B(_1852_),
    .Z(_1854_));
 XNOR2_X1 _5551_ (.A(_1842_),
    .B(_1843_),
    .ZN(_1855_));
 NAND2_X1 _5552_ (.A1(\section_1.yn2[6] ),
    .A2(\section_1.yn2[4] ),
    .ZN(_1856_));
 XOR2_X1 _5553_ (.A(\section_1.yn2[7] ),
    .B(\section_1.yn2[5] ),
    .Z(_1857_));
 XNOR2_X1 _5554_ (.A(_1652_),
    .B(_1857_),
    .ZN(_1859_));
 INV_X1 _5555_ (.A(_1859_),
    .ZN(_1860_));
 OAI22_X1 _5556_ (.A1(\section_1.yn2[5] ),
    .A2(_1652_),
    .B1(_1856_),
    .B2(_1860_),
    .ZN(_1861_));
 XNOR2_X1 _5557_ (.A(_0011_),
    .B(_1861_),
    .ZN(_1862_));
 XOR2_X1 _5558_ (.A(_1856_),
    .B(_1859_),
    .Z(_1863_));
 XNOR2_X1 _5559_ (.A(_1472_),
    .B(_1582_),
    .ZN(_1864_));
 XNOR2_X1 _5560_ (.A(_2717_),
    .B(_1864_),
    .ZN(_1865_));
 AOI22_X1 _5561_ (.A1(_0144_),
    .A2(_1864_),
    .B1(_1865_),
    .B2(\section_1.yn2[9] ),
    .ZN(_1866_));
 XOR2_X1 _5562_ (.A(_1585_),
    .B(_1586_),
    .Z(_1867_));
 XNOR2_X1 _5563_ (.A(_1866_),
    .B(_1867_),
    .ZN(_1868_));
 NAND2_X1 _5564_ (.A1(_0939_),
    .A2(_1868_),
    .ZN(_1870_));
 INV_X1 _5565_ (.A(_1867_),
    .ZN(_1871_));
 OAI21_X1 _5566_ (.A(_1870_),
    .B1(_1871_),
    .B2(_1866_),
    .ZN(_1872_));
 XOR2_X1 _5567_ (.A(_1823_),
    .B(_1824_),
    .Z(_1873_));
 XNOR2_X1 _5568_ (.A(_1872_),
    .B(_1873_),
    .ZN(_1874_));
 NOR2_X1 _5569_ (.A1(_1863_),
    .A2(_1874_),
    .ZN(_1875_));
 AOI21_X1 _5570_ (.A(_1875_),
    .B1(_1873_),
    .B2(_1872_),
    .ZN(_1876_));
 XNOR2_X1 _5571_ (.A(_1833_),
    .B(_1834_),
    .ZN(_1877_));
 XNOR2_X1 _5572_ (.A(_1876_),
    .B(_1877_),
    .ZN(_1878_));
 OR2_X1 _5573_ (.A1(_1862_),
    .A2(_1878_),
    .ZN(_1879_));
 OR2_X1 _5574_ (.A1(_1876_),
    .A2(_1877_),
    .ZN(_1881_));
 AOI21_X1 _5575_ (.A(_1855_),
    .B1(_1879_),
    .B2(_1881_),
    .ZN(_1882_));
 INV_X1 _5576_ (.A(_1882_),
    .ZN(_1883_));
 NAND3_X1 _5577_ (.A1(_1881_),
    .A2(_1879_),
    .A3(_1855_),
    .ZN(_1884_));
 NAND2_X1 _5578_ (.A1(_1883_),
    .A2(_1884_),
    .ZN(_1885_));
 NAND2_X1 _5579_ (.A1(_0011_),
    .A2(_1861_),
    .ZN(_1886_));
 OAI21_X1 _5580_ (.A(_1883_),
    .B1(_1885_),
    .B2(_1886_),
    .ZN(_1887_));
 XOR2_X1 _5581_ (.A(_1849_),
    .B(_1848_),
    .Z(_1888_));
 XNOR2_X1 _5582_ (.A(_1887_),
    .B(_1888_),
    .ZN(_1889_));
 XOR2_X1 _5583_ (.A(_0939_),
    .B(_1868_),
    .Z(_1890_));
 XNOR2_X1 _5584_ (.A(_1496_),
    .B(_1581_),
    .ZN(_1892_));
 AND2_X1 _5585_ (.A1(_2572_),
    .A2(_1892_),
    .ZN(_1893_));
 XNOR2_X1 _5586_ (.A(\section_1.yn2[9] ),
    .B(_1865_),
    .ZN(_1894_));
 XOR2_X1 _5587_ (.A(_1893_),
    .B(_1894_),
    .Z(_1895_));
 AND2_X1 _5588_ (.A1(_1830_),
    .A2(_1895_),
    .ZN(_1896_));
 NOR2_X1 _5589_ (.A1(_1893_),
    .A2(_1894_),
    .ZN(_1897_));
 OAI21_X1 _5590_ (.A(_1890_),
    .B1(_1896_),
    .B2(_1897_),
    .ZN(_1898_));
 NAND2_X1 _5591_ (.A1(\section_1.yn2[5] ),
    .A2(\section_1.yn2[3] ),
    .ZN(_1899_));
 XNOR2_X1 _5592_ (.A(\section_1.yn2[6] ),
    .B(\section_1.yn2[4] ),
    .ZN(_1900_));
 XOR2_X1 _5593_ (.A(_0938_),
    .B(_1900_),
    .Z(_1901_));
 XNOR2_X1 _5594_ (.A(_1899_),
    .B(_1901_),
    .ZN(_1903_));
 OR3_X1 _5595_ (.A1(_1897_),
    .A2(_1896_),
    .A3(_1890_),
    .ZN(_1904_));
 AND2_X1 _5596_ (.A1(_1898_),
    .A2(_1904_),
    .ZN(_1905_));
 NAND2_X1 _5597_ (.A1(_1903_),
    .A2(_1905_),
    .ZN(_1906_));
 NAND2_X1 _5598_ (.A1(_1898_),
    .A2(_1906_),
    .ZN(_1907_));
 XNOR2_X1 _5599_ (.A(_1863_),
    .B(_1874_),
    .ZN(_1908_));
 INV_X1 _5600_ (.A(_1908_),
    .ZN(_1909_));
 INV_X1 _5601_ (.A(_1901_),
    .ZN(_1910_));
 OAI22_X1 _5602_ (.A1(\section_1.yn2[4] ),
    .A2(_0938_),
    .B1(_1899_),
    .B2(_1910_),
    .ZN(_1911_));
 XOR2_X1 _5603_ (.A(_0012_),
    .B(_1911_),
    .Z(_1912_));
 XNOR2_X1 _5604_ (.A(_1907_),
    .B(_1908_),
    .ZN(_1914_));
 AOI22_X1 _5605_ (.A1(_1907_),
    .A2(_1909_),
    .B1(_1912_),
    .B2(_1914_),
    .ZN(_1915_));
 XNOR2_X1 _5606_ (.A(_1862_),
    .B(_1878_),
    .ZN(_1916_));
 NOR2_X1 _5607_ (.A1(_1915_),
    .A2(_1916_),
    .ZN(_1917_));
 XOR2_X1 _5608_ (.A(_1915_),
    .B(_1916_),
    .Z(_1918_));
 AND2_X1 _5609_ (.A1(_0012_),
    .A2(_1911_),
    .ZN(_1919_));
 AOI21_X1 _5610_ (.A(_1917_),
    .B1(_1918_),
    .B2(_1919_),
    .ZN(_1920_));
 XNOR2_X1 _5611_ (.A(_1886_),
    .B(_1885_),
    .ZN(_1921_));
 NOR2_X1 _5612_ (.A1(_1920_),
    .A2(_1921_),
    .ZN(_1922_));
 XOR2_X1 _5613_ (.A(_1920_),
    .B(_1921_),
    .Z(_1923_));
 XOR2_X1 _5614_ (.A(_0030_),
    .B(_1892_),
    .Z(_1925_));
 OR3_X1 _5615_ (.A1(_1514_),
    .A2(_1533_),
    .A3(_1579_),
    .ZN(_1926_));
 NAND2_X1 _5616_ (.A1(_1580_),
    .A2(_1926_),
    .ZN(_1927_));
 OR2_X1 _5617_ (.A1(_0008_),
    .A2(_1927_),
    .ZN(_1928_));
 XNOR2_X1 _5618_ (.A(_2504_),
    .B(_1927_),
    .ZN(_1929_));
 OR2_X1 _5619_ (.A1(_2443_),
    .A2(_1929_),
    .ZN(_1930_));
 AOI21_X1 _5620_ (.A(_1925_),
    .B1(_1928_),
    .B2(_1930_),
    .ZN(_1931_));
 XNOR2_X1 _5621_ (.A(\section_1.yn2[8] ),
    .B(\section_1.yn2[7] ),
    .ZN(_1932_));
 NAND2_X1 _5622_ (.A1(_1930_),
    .A2(_1928_),
    .ZN(_1933_));
 XOR2_X1 _5623_ (.A(_1933_),
    .B(_1925_),
    .Z(_1934_));
 NOR2_X1 _5624_ (.A1(_1932_),
    .A2(_1934_),
    .ZN(_1936_));
 OR2_X1 _5625_ (.A1(_1931_),
    .A2(_1936_),
    .ZN(_1937_));
 XOR2_X1 _5626_ (.A(_1830_),
    .B(_1895_),
    .Z(_1938_));
 NAND2_X1 _5627_ (.A1(\section_1.yn2[5] ),
    .A2(\section_1.yn2[4] ),
    .ZN(_1939_));
 NAND2_X1 _5628_ (.A1(\section_1.yn2[8] ),
    .A2(\section_1.yn2[7] ),
    .ZN(_1940_));
 XOR2_X1 _5629_ (.A(\section_1.yn2[5] ),
    .B(\section_1.yn2[3] ),
    .Z(_1941_));
 XNOR2_X1 _5630_ (.A(_1940_),
    .B(_1941_),
    .ZN(_1942_));
 XNOR2_X1 _5631_ (.A(_1939_),
    .B(_1942_),
    .ZN(_1943_));
 XOR2_X1 _5632_ (.A(_1937_),
    .B(_1938_),
    .Z(_1944_));
 AOI22_X1 _5633_ (.A1(_1937_),
    .A2(_1938_),
    .B1(_1943_),
    .B2(_1944_),
    .ZN(_1945_));
 XNOR2_X1 _5634_ (.A(_1903_),
    .B(_1905_),
    .ZN(_1947_));
 NOR2_X1 _5635_ (.A1(_1945_),
    .A2(_1947_),
    .ZN(_1948_));
 INV_X1 _5636_ (.A(_0013_),
    .ZN(_1949_));
 NAND3_X1 _5637_ (.A1(\section_1.yn2[8] ),
    .A2(\section_1.yn2[7] ),
    .A3(_1941_),
    .ZN(_1950_));
 NAND3_X1 _5638_ (.A1(\section_1.yn2[5] ),
    .A2(\section_1.yn2[4] ),
    .A3(_1942_),
    .ZN(_1951_));
 AND3_X1 _5639_ (.A1(_1949_),
    .A2(_1950_),
    .A3(_1951_),
    .ZN(_1952_));
 AOI21_X1 _5640_ (.A(_1949_),
    .B1(_1950_),
    .B2(_1951_),
    .ZN(_1953_));
 NOR2_X1 _5641_ (.A1(_1952_),
    .A2(_1953_),
    .ZN(_1954_));
 XOR2_X1 _5642_ (.A(_1945_),
    .B(_1947_),
    .Z(_1955_));
 AOI21_X1 _5643_ (.A(_1948_),
    .B1(_1954_),
    .B2(_1955_),
    .ZN(_1956_));
 XNOR2_X1 _5644_ (.A(_1912_),
    .B(_1914_),
    .ZN(_1958_));
 NOR2_X1 _5645_ (.A1(_1956_),
    .A2(_1958_),
    .ZN(_1959_));
 XOR2_X1 _5646_ (.A(_1956_),
    .B(_1958_),
    .Z(_1960_));
 AOI21_X1 _5647_ (.A(_1959_),
    .B1(_1960_),
    .B2(_1953_),
    .ZN(_1961_));
 XNOR2_X1 _5648_ (.A(_1919_),
    .B(_1918_),
    .ZN(_1962_));
 XOR2_X1 _5649_ (.A(_1961_),
    .B(_1962_),
    .Z(_1963_));
 XNOR2_X1 _5650_ (.A(_1576_),
    .B(_1578_),
    .ZN(_1964_));
 XNOR2_X1 _5651_ (.A(_2443_),
    .B(_1964_),
    .ZN(_1965_));
 OAI22_X1 _5652_ (.A1(_0001_),
    .A2(_1964_),
    .B1(_1965_),
    .B2(_2328_),
    .ZN(_1966_));
 XNOR2_X1 _5653_ (.A(\section_1.yn2[7] ),
    .B(_1929_),
    .ZN(_1967_));
 NAND2_X1 _5654_ (.A1(_1966_),
    .A2(_1967_),
    .ZN(_1969_));
 XNOR2_X1 _5655_ (.A(_1966_),
    .B(_1967_),
    .ZN(_1970_));
 OAI21_X1 _5656_ (.A(_1969_),
    .B1(_1970_),
    .B2(_1900_),
    .ZN(_1971_));
 XOR2_X1 _5657_ (.A(_1932_),
    .B(_1934_),
    .Z(_1972_));
 NAND2_X1 _5658_ (.A1(\section_1.yn2[3] ),
    .A2(\section_1.yn2[1] ),
    .ZN(_1973_));
 XOR2_X1 _5659_ (.A(\section_1.yn2[5] ),
    .B(\section_1.yn2[4] ),
    .Z(_1974_));
 XNOR2_X1 _5660_ (.A(_1856_),
    .B(_1974_),
    .ZN(_1975_));
 XNOR2_X1 _5661_ (.A(_1973_),
    .B(_1975_),
    .ZN(_1976_));
 XOR2_X1 _5662_ (.A(_1971_),
    .B(_1972_),
    .Z(_1977_));
 AOI22_X1 _5663_ (.A1(_1971_),
    .A2(_1972_),
    .B1(_1976_),
    .B2(_1977_),
    .ZN(_1978_));
 XNOR2_X1 _5664_ (.A(_1943_),
    .B(_1944_),
    .ZN(_1980_));
 NOR2_X1 _5665_ (.A1(_1978_),
    .A2(_1980_),
    .ZN(_1981_));
 NOR2_X1 _5666_ (.A1(_1528_),
    .A2(\section_1.yn2[0] ),
    .ZN(_1982_));
 NAND3_X1 _5667_ (.A1(\section_1.yn2[6] ),
    .A2(_2275_),
    .A3(\section_1.yn2[4] ),
    .ZN(_1983_));
 NAND3_X1 _5668_ (.A1(\section_1.yn2[3] ),
    .A2(\section_1.yn2[1] ),
    .A3(_1975_),
    .ZN(_1984_));
 NAND2_X1 _5669_ (.A1(_1983_),
    .A2(_1984_),
    .ZN(_1985_));
 XOR2_X1 _5670_ (.A(_0014_),
    .B(_1985_),
    .Z(_1986_));
 XOR2_X1 _5671_ (.A(_1982_),
    .B(_1986_),
    .Z(_1987_));
 XOR2_X1 _5672_ (.A(_1978_),
    .B(_1980_),
    .Z(_1988_));
 AOI21_X1 _5673_ (.A(_1981_),
    .B1(_1987_),
    .B2(_1988_),
    .ZN(_1989_));
 XNOR2_X1 _5674_ (.A(_1954_),
    .B(_1955_),
    .ZN(_1991_));
 NOR2_X1 _5675_ (.A1(_1989_),
    .A2(_1991_),
    .ZN(_1992_));
 NAND2_X1 _5676_ (.A1(_1982_),
    .A2(_1986_),
    .ZN(_1993_));
 OAI21_X1 _5677_ (.A(_1993_),
    .B1(_1983_),
    .B2(\section_1.yn2[1] ),
    .ZN(_1994_));
 XOR2_X1 _5678_ (.A(_1989_),
    .B(_1991_),
    .Z(_1995_));
 AOI21_X1 _5679_ (.A(_1992_),
    .B1(_1994_),
    .B2(_1995_),
    .ZN(_1996_));
 XNOR2_X1 _5680_ (.A(_1953_),
    .B(_1960_),
    .ZN(_1997_));
 NOR2_X1 _5681_ (.A1(_1996_),
    .A2(_1997_),
    .ZN(_1998_));
 XOR2_X1 _5682_ (.A(_1996_),
    .B(_1997_),
    .Z(_1999_));
 XOR2_X1 _5683_ (.A(_1987_),
    .B(_1988_),
    .Z(_2000_));
 XNOR2_X1 _5684_ (.A(\section_1.yn2[2] ),
    .B(\section_1.yn2[0] ),
    .ZN(_2002_));
 NAND2_X1 _5685_ (.A1(\section_1.yn2[2] ),
    .A2(\section_1.yn2[0] ),
    .ZN(_2003_));
 XNOR2_X1 _5686_ (.A(\section_1.yn2[3] ),
    .B(\section_1.yn2[1] ),
    .ZN(_2004_));
 XOR2_X1 _5687_ (.A(_1899_),
    .B(_2004_),
    .Z(_2005_));
 INV_X1 _5688_ (.A(_2005_),
    .ZN(_2006_));
 OAI22_X1 _5689_ (.A1(\section_1.yn2[1] ),
    .A2(_1899_),
    .B1(_2003_),
    .B2(_2006_),
    .ZN(_2007_));
 XNOR2_X1 _5690_ (.A(_2002_),
    .B(_2007_),
    .ZN(_2008_));
 XOR2_X1 _5691_ (.A(_1545_),
    .B(_1574_),
    .Z(_2009_));
 INV_X1 _5692_ (.A(_2009_),
    .ZN(_2010_));
 XNOR2_X1 _5693_ (.A(\section_1.yn2[6] ),
    .B(_2009_),
    .ZN(_2011_));
 OAI22_X1 _5694_ (.A1(_0003_),
    .A2(_2010_),
    .B1(_2011_),
    .B2(_2275_),
    .ZN(_2013_));
 INV_X1 _5695_ (.A(_2013_),
    .ZN(_2014_));
 XNOR2_X1 _5696_ (.A(_2328_),
    .B(_1965_),
    .ZN(_2015_));
 OR2_X1 _5697_ (.A1(_2014_),
    .A2(_2015_),
    .ZN(_2016_));
 XNOR2_X1 _5698_ (.A(_2014_),
    .B(_2015_),
    .ZN(_2017_));
 INV_X1 _5699_ (.A(_1941_),
    .ZN(_2018_));
 OAI21_X1 _5700_ (.A(_2016_),
    .B1(_2017_),
    .B2(_2018_),
    .ZN(_2019_));
 XOR2_X1 _5701_ (.A(_1900_),
    .B(_1970_),
    .Z(_2020_));
 XOR2_X1 _5702_ (.A(_2019_),
    .B(_2020_),
    .Z(_2021_));
 XNOR2_X1 _5703_ (.A(_2003_),
    .B(_2005_),
    .ZN(_2022_));
 AOI22_X1 _5704_ (.A1(_2019_),
    .A2(_2020_),
    .B1(_2021_),
    .B2(_2022_),
    .ZN(_2024_));
 XNOR2_X1 _5705_ (.A(_1976_),
    .B(_1977_),
    .ZN(_2025_));
 XOR2_X1 _5706_ (.A(_2024_),
    .B(_2025_),
    .Z(_2026_));
 INV_X1 _5707_ (.A(_2026_),
    .ZN(_2027_));
 NOR2_X1 _5708_ (.A1(_2008_),
    .A2(_2027_),
    .ZN(_2028_));
 NOR2_X1 _5709_ (.A1(_2024_),
    .A2(_2025_),
    .ZN(_2029_));
 OAI21_X1 _5710_ (.A(_2000_),
    .B1(_2028_),
    .B2(_2029_),
    .ZN(_2030_));
 INV_X1 _5711_ (.A(_2030_),
    .ZN(_2031_));
 NOR2_X1 _5712_ (.A1(_2029_),
    .A2(_2028_),
    .ZN(_2032_));
 XNOR2_X1 _5713_ (.A(_2032_),
    .B(_2000_),
    .ZN(_2033_));
 NAND2_X1 _5714_ (.A1(_2002_),
    .A2(_2007_),
    .ZN(_2035_));
 INV_X1 _5715_ (.A(_2035_),
    .ZN(_2036_));
 AOI21_X1 _5716_ (.A(_2031_),
    .B1(_2033_),
    .B2(_2036_),
    .ZN(_2037_));
 XNOR2_X1 _5717_ (.A(_1994_),
    .B(_1995_),
    .ZN(_2038_));
 XOR2_X1 _5718_ (.A(_2037_),
    .B(_2038_),
    .Z(_2039_));
 XNOR2_X1 _5719_ (.A(_2021_),
    .B(_2022_),
    .ZN(_2040_));
 XNOR2_X1 _5720_ (.A(_1941_),
    .B(_2017_),
    .ZN(_2041_));
 XNOR2_X1 _5721_ (.A(_1571_),
    .B(_1573_),
    .ZN(_2042_));
 XNOR2_X1 _5722_ (.A(_2275_),
    .B(_2042_),
    .ZN(_2043_));
 OAI22_X1 _5723_ (.A1(_0009_),
    .A2(_2042_),
    .B1(_2043_),
    .B2(_0916_),
    .ZN(_2044_));
 INV_X1 _5724_ (.A(_2044_),
    .ZN(_2046_));
 XNOR2_X1 _5725_ (.A(_2275_),
    .B(_2011_),
    .ZN(_2047_));
 XNOR2_X1 _5726_ (.A(_2046_),
    .B(_2047_),
    .ZN(_2048_));
 XNOR2_X1 _5727_ (.A(\section_1.yn2[4] ),
    .B(\section_1.yn2[2] ),
    .ZN(_2049_));
 NOR2_X1 _5728_ (.A1(_2048_),
    .A2(_2049_),
    .ZN(_2050_));
 NOR2_X1 _5729_ (.A1(_2046_),
    .A2(_2047_),
    .ZN(_2051_));
 OAI21_X1 _5730_ (.A(_2041_),
    .B1(_2050_),
    .B2(_2051_),
    .ZN(_2052_));
 OR3_X1 _5731_ (.A1(_2051_),
    .A2(_2050_),
    .A3(_2041_),
    .ZN(_2053_));
 AND2_X1 _5732_ (.A1(_2052_),
    .A2(_2053_),
    .ZN(_2054_));
 NAND2_X1 _5733_ (.A1(\section_1.yn2[4] ),
    .A2(\section_1.yn2[2] ),
    .ZN(_2055_));
 XOR2_X1 _5734_ (.A(_2002_),
    .B(_2055_),
    .Z(_2057_));
 NAND2_X1 _5735_ (.A1(_2054_),
    .A2(_2057_),
    .ZN(_2058_));
 AOI21_X1 _5736_ (.A(_2040_),
    .B1(_2058_),
    .B2(_2052_),
    .ZN(_2059_));
 AND3_X1 _5737_ (.A1(_2052_),
    .A2(_2058_),
    .A3(_2040_),
    .ZN(_2060_));
 NOR2_X1 _5738_ (.A1(_2059_),
    .A2(_2060_),
    .ZN(_2061_));
 NOR2_X1 _5739_ (.A1(\section_1.yn2[0] ),
    .A2(_2055_),
    .ZN(_2062_));
 AOI21_X1 _5740_ (.A(_2059_),
    .B1(_2061_),
    .B2(_2062_),
    .ZN(_2063_));
 XOR2_X1 _5741_ (.A(_2008_),
    .B(_2026_),
    .Z(_2064_));
 NOR2_X1 _5742_ (.A1(_2063_),
    .A2(_2064_),
    .ZN(_2065_));
 XNOR2_X1 _5743_ (.A(_2035_),
    .B(_2033_),
    .ZN(_2066_));
 AND2_X1 _5744_ (.A1(_2065_),
    .A2(_2066_),
    .ZN(_2068_));
 XNOR2_X1 _5745_ (.A(_2065_),
    .B(_2066_),
    .ZN(_2069_));
 XOR2_X1 _5746_ (.A(_2062_),
    .B(_2061_),
    .Z(_2070_));
 XNOR2_X1 _5747_ (.A(_1568_),
    .B(_1570_),
    .ZN(_2071_));
 XNOR2_X1 _5748_ (.A(_0916_),
    .B(_2071_),
    .ZN(_2072_));
 OAI22_X1 _5749_ (.A1(_0011_),
    .A2(_2071_),
    .B1(_2072_),
    .B2(_0917_),
    .ZN(_2073_));
 XNOR2_X1 _5750_ (.A(\section_1.yn2[4] ),
    .B(_2043_),
    .ZN(_2074_));
 NAND2_X1 _5751_ (.A1(_2073_),
    .A2(_2074_),
    .ZN(_2075_));
 XNOR2_X1 _5752_ (.A(_2073_),
    .B(_2074_),
    .ZN(_2076_));
 OAI21_X1 _5753_ (.A(_2075_),
    .B1(_2076_),
    .B2(_2004_),
    .ZN(_2077_));
 XOR2_X1 _5754_ (.A(_2048_),
    .B(_2049_),
    .Z(_2079_));
 NAND2_X1 _5755_ (.A1(_2077_),
    .A2(_2079_),
    .ZN(_2080_));
 XNOR2_X1 _5756_ (.A(_2077_),
    .B(_2079_),
    .ZN(_2081_));
 NAND2_X1 _5757_ (.A1(_0917_),
    .A2(\section_1.yn2[1] ),
    .ZN(_2082_));
 OAI21_X1 _5758_ (.A(_2080_),
    .B1(_2081_),
    .B2(_2082_),
    .ZN(_2083_));
 INV_X1 _5759_ (.A(_2083_),
    .ZN(_2084_));
 XNOR2_X1 _5760_ (.A(_2054_),
    .B(_2057_),
    .ZN(_2085_));
 XNOR2_X1 _5761_ (.A(_2084_),
    .B(_2085_),
    .ZN(_2086_));
 NOR2_X1 _5762_ (.A1(_1973_),
    .A2(_2086_),
    .ZN(_2087_));
 NOR2_X1 _5763_ (.A1(_2084_),
    .A2(_2085_),
    .ZN(_2088_));
 OAI21_X1 _5764_ (.A(_2070_),
    .B1(_2087_),
    .B2(_2088_),
    .ZN(_2090_));
 XOR2_X1 _5765_ (.A(_2063_),
    .B(_2064_),
    .Z(_2091_));
 XNOR2_X1 _5766_ (.A(_2090_),
    .B(_2091_),
    .ZN(_2092_));
 OR3_X1 _5767_ (.A1(_2088_),
    .A2(_2087_),
    .A3(_2070_),
    .ZN(_2093_));
 AND2_X1 _5768_ (.A1(_2090_),
    .A2(_2093_),
    .ZN(_2094_));
 NAND2_X1 _5769_ (.A1(_1528_),
    .A2(\section_1.yn2[0] ),
    .ZN(_2095_));
 XNOR2_X1 _5770_ (.A(_1566_),
    .B(_1567_),
    .ZN(_2096_));
 XNOR2_X1 _5771_ (.A(_0917_),
    .B(_2096_),
    .ZN(_2097_));
 OAI22_X1 _5772_ (.A1(_0012_),
    .A2(_2096_),
    .B1(_2097_),
    .B2(_1528_),
    .ZN(_2098_));
 XNOR2_X1 _5773_ (.A(\section_1.yn2[3] ),
    .B(_2072_),
    .ZN(_2099_));
 NAND2_X1 _5774_ (.A1(_2098_),
    .A2(_2099_),
    .ZN(_2101_));
 XNOR2_X1 _5775_ (.A(_2098_),
    .B(_2099_),
    .ZN(_2102_));
 OAI21_X1 _5776_ (.A(_2101_),
    .B1(_2102_),
    .B2(_2002_),
    .ZN(_2103_));
 XOR2_X1 _5777_ (.A(_2004_),
    .B(_2076_),
    .Z(_2104_));
 XNOR2_X1 _5778_ (.A(_2103_),
    .B(_2104_),
    .ZN(_2105_));
 NOR2_X1 _5779_ (.A1(_2095_),
    .A2(_2105_),
    .ZN(_2106_));
 AOI21_X1 _5780_ (.A(_2106_),
    .B1(_2104_),
    .B2(_2103_),
    .ZN(_2107_));
 XNOR2_X1 _5781_ (.A(_2081_),
    .B(_2082_),
    .ZN(_2108_));
 XNOR2_X1 _5782_ (.A(_2107_),
    .B(_2108_),
    .ZN(_2109_));
 OR2_X1 _5783_ (.A1(_2003_),
    .A2(_2109_),
    .ZN(_2110_));
 OAI21_X1 _5784_ (.A(_2110_),
    .B1(_2108_),
    .B2(_2107_),
    .ZN(_2112_));
 XOR2_X1 _5785_ (.A(_1973_),
    .B(_2086_),
    .Z(_2113_));
 NOR2_X1 _5786_ (.A1(_2112_),
    .A2(_2113_),
    .ZN(_2114_));
 NAND2_X1 _5787_ (.A1(_2003_),
    .A2(_2109_),
    .ZN(_2115_));
 XNOR2_X1 _5788_ (.A(_1563_),
    .B(_1565_),
    .ZN(_2116_));
 XNOR2_X1 _5789_ (.A(_1528_),
    .B(_2116_),
    .ZN(_2117_));
 OAI22_X1 _5790_ (.A1(_0013_),
    .A2(_2116_),
    .B1(_2117_),
    .B2(_1330_),
    .ZN(_2118_));
 XNOR2_X1 _5791_ (.A(\section_1.yn2[2] ),
    .B(_2097_),
    .ZN(_2119_));
 NAND2_X1 _5792_ (.A1(_2118_),
    .A2(_2119_),
    .ZN(_2120_));
 XNOR2_X1 _5793_ (.A(_2118_),
    .B(_2119_),
    .ZN(_2121_));
 OR2_X1 _5794_ (.A1(_1330_),
    .A2(_2121_),
    .ZN(_2123_));
 XNOR2_X1 _5795_ (.A(_2002_),
    .B(_2102_),
    .ZN(_2124_));
 NAND3_X1 _5796_ (.A1(_2120_),
    .A2(_2123_),
    .A3(_2124_),
    .ZN(_2125_));
 AOI21_X1 _5797_ (.A(_2124_),
    .B1(_2123_),
    .B2(_2120_),
    .ZN(_2126_));
 XNOR2_X1 _5798_ (.A(\section_1.yn2[1] ),
    .B(_2121_),
    .ZN(_2127_));
 XNOR2_X1 _5799_ (.A(_1560_),
    .B(_1562_),
    .ZN(_2128_));
 XNOR2_X1 _5800_ (.A(_1330_),
    .B(_2128_),
    .ZN(_2129_));
 OAI22_X1 _5801_ (.A1(_0014_),
    .A2(_2128_),
    .B1(_2129_),
    .B2(_2386_),
    .ZN(_2130_));
 XNOR2_X1 _5802_ (.A(\section_1.yn2[1] ),
    .B(_2117_),
    .ZN(_2131_));
 XOR2_X1 _5803_ (.A(_2130_),
    .B(_2131_),
    .Z(_2132_));
 AND2_X1 _5804_ (.A1(\section_1.yn2[0] ),
    .A2(_2132_),
    .ZN(_2134_));
 AND2_X1 _5805_ (.A1(_2130_),
    .A2(_2131_),
    .ZN(_2135_));
 OAI21_X1 _5806_ (.A(_2127_),
    .B1(_2134_),
    .B2(_2135_),
    .ZN(_2136_));
 NOR3_X1 _5807_ (.A1(_2135_),
    .A2(_2134_),
    .A3(_2127_),
    .ZN(_2137_));
 AOI21_X1 _5808_ (.A(_1559_),
    .B1(\section_1.t1[0] ),
    .B2(\coll_reg[0] ),
    .ZN(_2138_));
 INV_X1 _5809_ (.A(_0015_),
    .ZN(_2139_));
 NAND2_X1 _5810_ (.A1(_2139_),
    .A2(_1560_),
    .ZN(_2140_));
 NAND2_X1 _5811_ (.A1(_2386_),
    .A2(_2129_),
    .ZN(_2141_));
 OAI21_X1 _5812_ (.A(_2141_),
    .B1(_2132_),
    .B2(_2129_),
    .ZN(_2142_));
 OR4_X1 _5813_ (.A1(_2134_),
    .A2(_2138_),
    .A3(_2140_),
    .A4(_2142_),
    .ZN(_2143_));
 OAI21_X1 _5814_ (.A(_2136_),
    .B1(_2137_),
    .B2(_2143_),
    .ZN(_2145_));
 OAI221_X1 _5815_ (.A(_2125_),
    .B1(_2126_),
    .B2(_2145_),
    .C1(_2105_),
    .C2(_2095_),
    .ZN(_2146_));
 AOI21_X1 _5816_ (.A(_2146_),
    .B1(_2105_),
    .B2(_2095_),
    .ZN(_2147_));
 NAND3_X1 _5817_ (.A1(_2110_),
    .A2(_2115_),
    .A3(_2147_),
    .ZN(_2148_));
 NOR2_X1 _5818_ (.A1(_2114_),
    .A2(_2148_),
    .ZN(_2149_));
 AND2_X1 _5819_ (.A1(_2112_),
    .A2(_2113_),
    .ZN(_2150_));
 OAI211_X1 _5820_ (.A(_2092_),
    .B(_2094_),
    .C1(_2149_),
    .C2(_2150_),
    .ZN(_2151_));
 INV_X1 _5821_ (.A(_2091_),
    .ZN(_2152_));
 OAI21_X1 _5822_ (.A(_2151_),
    .B1(_2152_),
    .B2(_2090_),
    .ZN(_2153_));
 INV_X1 _5823_ (.A(_2153_),
    .ZN(_2154_));
 NOR2_X1 _5824_ (.A1(_2069_),
    .A2(_2154_),
    .ZN(_2156_));
 OAI21_X1 _5825_ (.A(_2039_),
    .B1(_2068_),
    .B2(_2156_),
    .ZN(_2157_));
 OAI21_X1 _5826_ (.A(_2157_),
    .B1(_2038_),
    .B2(_2037_),
    .ZN(_2158_));
 AND2_X1 _5827_ (.A1(_1999_),
    .A2(_2158_),
    .ZN(_2159_));
 OAI21_X1 _5828_ (.A(_1963_),
    .B1(_1998_),
    .B2(_2159_),
    .ZN(_2160_));
 OAI21_X1 _5829_ (.A(_2160_),
    .B1(_1962_),
    .B2(_1961_),
    .ZN(_2161_));
 AOI21_X1 _5830_ (.A(_1922_),
    .B1(_1923_),
    .B2(_2161_),
    .ZN(_2162_));
 NOR2_X1 _5831_ (.A1(_1889_),
    .A2(_2162_),
    .ZN(_2163_));
 AND2_X1 _5832_ (.A1(_1887_),
    .A2(_1888_),
    .ZN(_2164_));
 OAI21_X1 _5833_ (.A(_1854_),
    .B1(_2163_),
    .B2(_2164_),
    .ZN(_2165_));
 AND2_X1 _5834_ (.A1(_1853_),
    .A2(_2165_),
    .ZN(_2167_));
 OAI21_X1 _5835_ (.A(_1818_),
    .B1(_1819_),
    .B2(_2167_),
    .ZN(_2168_));
 OAI21_X1 _5836_ (.A(_1813_),
    .B1(_1816_),
    .B2(_1766_),
    .ZN(_2169_));
 NAND2_X1 _5837_ (.A1(_0008_),
    .A2(_1767_),
    .ZN(_2170_));
 NAND2_X1 _5838_ (.A1(\section_1.yn2[9] ),
    .A2(_2717_),
    .ZN(_2171_));
 NOR3_X1 _5839_ (.A1(\section_1.yn2[9] ),
    .A2(_2717_),
    .A3(_1807_),
    .ZN(_2172_));
 AOI21_X1 _5840_ (.A(_2172_),
    .B1(_1806_),
    .B2(_1774_),
    .ZN(_2173_));
 XNOR2_X1 _5841_ (.A(_1654_),
    .B(_1805_),
    .ZN(_2174_));
 NAND2_X1 _5842_ (.A1(_0144_),
    .A2(_2174_),
    .ZN(_2175_));
 NAND2_X1 _5843_ (.A1(_1777_),
    .A2(_1800_),
    .ZN(_2176_));
 NAND2_X1 _5844_ (.A1(_2176_),
    .A2(_1804_),
    .ZN(_2178_));
 NOR2_X1 _5845_ (.A1(_1780_),
    .A2(_1798_),
    .ZN(_2179_));
 AOI21_X1 _5846_ (.A(_2179_),
    .B1(_1799_),
    .B2(_1778_),
    .ZN(_2180_));
 NOR3_X1 _5847_ (.A1(_2452_),
    .A2(_2588_),
    .A3(_1782_),
    .ZN(_2181_));
 NAND2_X1 _5848_ (.A1(_1786_),
    .A2(_1796_),
    .ZN(_2182_));
 OAI21_X1 _5849_ (.A(_2182_),
    .B1(_1797_),
    .B2(_1785_),
    .ZN(_2183_));
 AOI21_X1 _5850_ (.A(_2659_),
    .B1(_1404_),
    .B2(\coll_reg[9] ),
    .ZN(_2184_));
 NAND2_X1 _5851_ (.A1(_1789_),
    .A2(_1794_),
    .ZN(_2185_));
 OAI211_X1 _5852_ (.A(_1285_),
    .B(_0010_),
    .C1(_0927_),
    .C2(\in_reg1[10] ),
    .ZN(_2186_));
 INV_X1 _5853_ (.A(_1787_),
    .ZN(_2187_));
 OAI211_X1 _5854_ (.A(_2185_),
    .B(_2186_),
    .C1(_1795_),
    .C2(_2187_),
    .ZN(_2189_));
 XOR2_X1 _5855_ (.A(_2184_),
    .B(_2189_),
    .Z(_2190_));
 XOR2_X1 _5856_ (.A(_2183_),
    .B(_2190_),
    .Z(_2191_));
 XOR2_X1 _5857_ (.A(_2181_),
    .B(_2191_),
    .Z(_2192_));
 XNOR2_X1 _5858_ (.A(_2180_),
    .B(_2192_),
    .ZN(_2193_));
 XOR2_X1 _5859_ (.A(_2178_),
    .B(_2193_),
    .Z(_2194_));
 XNOR2_X1 _5860_ (.A(\section_1.yn2[10] ),
    .B(_2194_),
    .ZN(_2195_));
 XNOR2_X1 _5861_ (.A(_2175_),
    .B(_2195_),
    .ZN(_2196_));
 XNOR2_X1 _5862_ (.A(_2173_),
    .B(_2196_),
    .ZN(_2197_));
 XNOR2_X1 _5863_ (.A(_2171_),
    .B(_2197_),
    .ZN(_2198_));
 AND2_X1 _5864_ (.A1(_1768_),
    .A2(_1809_),
    .ZN(_2200_));
 AND2_X1 _5865_ (.A1(_1771_),
    .A2(_1808_),
    .ZN(_2201_));
 OAI21_X1 _5866_ (.A(_2198_),
    .B1(_2200_),
    .B2(_2201_),
    .ZN(_2202_));
 OR3_X1 _5867_ (.A1(_2201_),
    .A2(_2200_),
    .A3(_2198_),
    .ZN(_2203_));
 AND2_X1 _5868_ (.A1(_2202_),
    .A2(_2203_),
    .ZN(_2204_));
 XNOR2_X1 _5869_ (.A(_2170_),
    .B(_2204_),
    .ZN(_2205_));
 XOR2_X1 _5870_ (.A(_2169_),
    .B(_2205_),
    .Z(_2206_));
 XOR2_X1 _5871_ (.A(_2168_),
    .B(_2206_),
    .Z(_2207_));
 XOR2_X1 _5872_ (.A(_1764_),
    .B(_1817_),
    .Z(_2208_));
 XNOR2_X1 _5873_ (.A(_2208_),
    .B(_2167_),
    .ZN(_2209_));
 OR3_X1 _5874_ (.A1(_2164_),
    .A2(_2163_),
    .A3(_1854_),
    .ZN(_2211_));
 AND2_X1 _5875_ (.A1(_2165_),
    .A2(_2211_),
    .ZN(_2212_));
 XOR2_X1 _5876_ (.A(_1889_),
    .B(_2162_),
    .Z(_2213_));
 XOR2_X1 _5877_ (.A(_1923_),
    .B(_2161_),
    .Z(_2214_));
 OR3_X1 _5878_ (.A1(_1963_),
    .A2(_1998_),
    .A3(_2159_),
    .ZN(_2215_));
 AND2_X1 _5879_ (.A1(_2160_),
    .A2(_2215_),
    .ZN(_2216_));
 OR3_X1 _5880_ (.A1(_2039_),
    .A2(_2068_),
    .A3(_2156_),
    .ZN(_2217_));
 AND2_X1 _5881_ (.A1(_2157_),
    .A2(_2217_),
    .ZN(_2218_));
 XNOR2_X1 _5882_ (.A(_2150_),
    .B(_2094_),
    .ZN(_2219_));
 XNOR2_X1 _5883_ (.A(_2149_),
    .B(_2219_),
    .ZN(_2220_));
 OAI21_X1 _5884_ (.A(_2094_),
    .B1(_2149_),
    .B2(_2150_),
    .ZN(_2222_));
 XNOR2_X1 _5885_ (.A(_2092_),
    .B(_2222_),
    .ZN(_2223_));
 AND2_X1 _5886_ (.A1(_2220_),
    .A2(_2223_),
    .ZN(_2224_));
 XNOR2_X1 _5887_ (.A(_2069_),
    .B(_2153_),
    .ZN(_2225_));
 AND2_X1 _5888_ (.A1(_2224_),
    .A2(_2225_),
    .ZN(_2226_));
 AND2_X1 _5889_ (.A1(_2218_),
    .A2(_2226_),
    .ZN(_2227_));
 XOR2_X1 _5890_ (.A(_1999_),
    .B(_2158_),
    .Z(_2228_));
 AND2_X1 _5891_ (.A1(_2227_),
    .A2(_2228_),
    .ZN(_2229_));
 AND2_X1 _5892_ (.A1(_2216_),
    .A2(_2229_),
    .ZN(_2230_));
 AND2_X1 _5893_ (.A1(_2214_),
    .A2(_2230_),
    .ZN(_2231_));
 AND2_X1 _5894_ (.A1(_2213_),
    .A2(_2231_),
    .ZN(_2233_));
 AND2_X1 _5895_ (.A1(_2212_),
    .A2(_2233_),
    .ZN(_2234_));
 AND2_X1 _5896_ (.A1(_2209_),
    .A2(_2234_),
    .ZN(_2235_));
 OAI21_X1 _5897_ (.A(_1253_),
    .B1(_2207_),
    .B2(_2235_),
    .ZN(_2236_));
 AOI21_X1 _5898_ (.A(_2236_),
    .B1(_2235_),
    .B2(_2207_),
    .ZN(_0042_));
 NOR2_X1 _5899_ (.A1(_2209_),
    .A2(_2234_),
    .ZN(_2237_));
 NOR3_X1 _5900_ (.A1(rst),
    .A2(_2235_),
    .A3(_2237_),
    .ZN(_0041_));
 NOR2_X1 _5901_ (.A1(_2212_),
    .A2(_2233_),
    .ZN(_2238_));
 NOR3_X1 _5902_ (.A1(rst),
    .A2(_2234_),
    .A3(_2238_),
    .ZN(_0040_));
 NOR2_X1 _5903_ (.A1(_2213_),
    .A2(_2231_),
    .ZN(_2239_));
 NOR3_X1 _5904_ (.A1(rst),
    .A2(_2233_),
    .A3(_2239_),
    .ZN(_0039_));
 NOR2_X1 _5905_ (.A1(_2214_),
    .A2(_2230_),
    .ZN(_2241_));
 NOR3_X1 _5906_ (.A1(rst),
    .A2(_2231_),
    .A3(_2241_),
    .ZN(_0038_));
 NOR2_X1 _5907_ (.A1(_2216_),
    .A2(_2229_),
    .ZN(_2242_));
 NOR3_X1 _5908_ (.A1(rst),
    .A2(_2230_),
    .A3(_2242_),
    .ZN(_0037_));
 NOR2_X1 _5909_ (.A1(_2227_),
    .A2(_2228_),
    .ZN(_2243_));
 NOR3_X1 _5910_ (.A1(rst),
    .A2(_2229_),
    .A3(_2243_),
    .ZN(_0036_));
 NOR2_X1 _5911_ (.A1(_2218_),
    .A2(_2226_),
    .ZN(_2244_));
 NOR3_X1 _5912_ (.A1(rst),
    .A2(_2227_),
    .A3(_2244_),
    .ZN(_0035_));
 NOR2_X1 _5913_ (.A1(_2224_),
    .A2(_2225_),
    .ZN(_2245_));
 NOR3_X1 _5914_ (.A1(rst),
    .A2(_2226_),
    .A3(_2245_),
    .ZN(_0034_));
 NAND2_X1 _5915_ (.A1(_2207_),
    .A2(_2235_),
    .ZN(_2247_));
 AND2_X1 _5916_ (.A1(_2169_),
    .A2(_2205_),
    .ZN(_2248_));
 AOI21_X1 _5917_ (.A(_2248_),
    .B1(_2206_),
    .B2(_2168_),
    .ZN(_2249_));
 NAND3_X1 _5918_ (.A1(_0008_),
    .A2(_1767_),
    .A3(_2204_),
    .ZN(_2250_));
 NAND2_X1 _5919_ (.A1(_2202_),
    .A2(_2250_),
    .ZN(_2251_));
 INV_X1 _5920_ (.A(_2197_),
    .ZN(_2252_));
 NAND2_X1 _5921_ (.A1(_2171_),
    .A2(_2252_),
    .ZN(_2253_));
 OAI21_X1 _5922_ (.A(_2253_),
    .B1(_2196_),
    .B2(_2173_),
    .ZN(_2254_));
 NOR3_X1 _5923_ (.A1(_0004_),
    .A2(_2174_),
    .A3(_2195_),
    .ZN(_2255_));
 NAND3_X1 _5924_ (.A1(\section_1.yn2[9] ),
    .A2(\section_1.yn2[10] ),
    .A3(_0030_),
    .ZN(_2257_));
 INV_X1 _5925_ (.A(_2192_),
    .ZN(_2258_));
 NOR2_X1 _5926_ (.A1(_2180_),
    .A2(_2258_),
    .ZN(_2259_));
 AOI21_X1 _5927_ (.A(_2259_),
    .B1(_2193_),
    .B2(_2178_),
    .ZN(_2260_));
 AOI22_X1 _5928_ (.A1(_2183_),
    .A2(_2190_),
    .B1(_2191_),
    .B2(_2181_),
    .ZN(_2261_));
 AOI211_X1 _5929_ (.A(_2659_),
    .B(_2189_),
    .C1(_1404_),
    .C2(\coll_reg[9] ),
    .ZN(_2262_));
 XNOR2_X1 _5930_ (.A(_2661_),
    .B(_2262_),
    .ZN(_2263_));
 XNOR2_X1 _5931_ (.A(_2261_),
    .B(_2263_),
    .ZN(_2264_));
 XNOR2_X1 _5932_ (.A(_2260_),
    .B(_2264_),
    .ZN(_2265_));
 XNOR2_X1 _5933_ (.A(_2257_),
    .B(_2265_),
    .ZN(_2266_));
 XOR2_X1 _5934_ (.A(_2255_),
    .B(_2266_),
    .Z(_2268_));
 XNOR2_X1 _5935_ (.A(_2254_),
    .B(_2268_),
    .ZN(_2269_));
 XNOR2_X1 _5936_ (.A(_2251_),
    .B(_2269_),
    .ZN(_2270_));
 XNOR2_X1 _5937_ (.A(_2249_),
    .B(_2270_),
    .ZN(_2271_));
 OAI21_X1 _5938_ (.A(_1253_),
    .B1(_2247_),
    .B2(_2271_),
    .ZN(_2272_));
 AOI21_X1 _5939_ (.A(_2272_),
    .B1(_2271_),
    .B2(_2247_),
    .ZN(_0033_));
 NOR2_X1 _5940_ (.A1(_2220_),
    .A2(_2223_),
    .ZN(_2273_));
 NOR3_X1 _5941_ (.A1(rst),
    .A2(_2224_),
    .A3(_2273_),
    .ZN(_0032_));
 DFF_X1 \coll_reg[0]$_SDFF_PP0_  (.D(_0032_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\coll_reg[0] ),
    .QN(_3014_));
 DFF_X1 \coll_reg[10]$_SDFF_PP0_  (.D(_0033_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\coll_reg[10] ),
    .QN(_0006_));
 DFF_X1 \coll_reg[1]$_SDFF_PP0_  (.D(_0034_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\coll_reg[1] ),
    .QN(_3013_));
 DFF_X1 \coll_reg[2]$_SDFF_PP0_  (.D(_0035_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\coll_reg[2] ),
    .QN(_3012_));
 DFF_X1 \coll_reg[3]$_SDFF_PP0_  (.D(_0036_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\coll_reg[3] ),
    .QN(_3011_));
 DFF_X1 \coll_reg[4]$_SDFF_PP0_  (.D(_0037_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\coll_reg[4] ),
    .QN(_3010_));
 DFF_X1 \coll_reg[5]$_SDFF_PP0_  (.D(_0038_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\coll_reg[5] ),
    .QN(_0007_));
 DFF_X1 \coll_reg[6]$_SDFF_PP0_  (.D(_0039_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\coll_reg[6] ),
    .QN(_3009_));
 DFF_X1 \coll_reg[7]$_SDFF_PP0_  (.D(_0040_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\coll_reg[7] ),
    .QN(_3008_));
 DFF_X1 \coll_reg[8]$_SDFF_PP0_  (.D(_0041_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\coll_reg[8] ),
    .QN(_0005_));
 DFF_X1 \coll_reg[9]$_SDFF_PP0_  (.D(_0042_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\coll_reg[9] ),
    .QN(_0000_));
 DFF_X1 \in_reg1[0]$_SDFF_PP0_  (.D(_0043_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\in_reg1[0] ),
    .QN(_3007_));
 DFF_X1 \in_reg1[10]$_SDFF_PP0_  (.D(_0044_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\in_reg1[10] ),
    .QN(_0010_));
 DFF_X1 \in_reg1[1]$_SDFF_PP0_  (.D(_0045_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\in_reg1[1] ),
    .QN(_3006_));
 DFF_X1 \in_reg1[2]$_SDFF_PP0_  (.D(_0046_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\in_reg1[2] ),
    .QN(_3005_));
 DFF_X1 \in_reg1[3]$_SDFF_PP0_  (.D(_0047_),
    .CK(clknet_3_7__leaf_clk),
    .Q(\in_reg1[3] ),
    .QN(_3004_));
 DFF_X1 \in_reg1[4]$_SDFF_PP0_  (.D(_0048_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\in_reg1[4] ),
    .QN(_3003_));
 DFF_X1 \in_reg1[5]$_SDFF_PP0_  (.D(_0049_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\in_reg1[5] ),
    .QN(_3002_));
 DFF_X1 \in_reg1[6]$_SDFF_PP0_  (.D(_0050_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\in_reg1[6] ),
    .QN(_3001_));
 DFF_X1 \in_reg1[7]$_SDFF_PP0_  (.D(_0051_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\in_reg1[7] ),
    .QN(_3000_));
 DFF_X1 \in_reg1[8]$_SDFF_PP0_  (.D(_0052_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\in_reg1[8] ),
    .QN(_2999_));
 DFF_X1 \in_reg1[9]$_SDFF_PP0_  (.D(_0053_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\in_reg1[9] ),
    .QN(_2998_));
 DFF_X1 \section_1.t1[0]$_SDFF_PP0_  (.D(net30),
    .CK(clknet_3_0__leaf_clk),
    .Q(\section_1.t1[0] ),
    .QN(_2997_));
 DFF_X1 \section_1.t1[1]$_SDFF_PP0_  (.D(_0055_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\section_1.t1[1] ),
    .QN(_2996_));
 DFF_X1 \section_1.t1[2]$_SDFF_PP0_  (.D(_0056_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\section_1.t1[2] ),
    .QN(_2995_));
 DFF_X1 \section_1.t1[3]$_SDFF_PP0_  (.D(_0057_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\section_1.t1[3] ),
    .QN(_2994_));
 DFF_X1 \section_1.t1[4]$_SDFF_PP0_  (.D(_0058_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\section_1.t1[4] ),
    .QN(_2993_));
 DFF_X1 \section_1.xn1[10]$_SDFF_PP0_  (.D(net16),
    .CK(clknet_3_2__leaf_clk),
    .Q(\section_1.xn1[10] ),
    .QN(_2992_));
 DFF_X1 \section_1.xn1[5]$_SDFF_PP0_  (.D(net19),
    .CK(clknet_3_0__leaf_clk),
    .Q(\section_1.xn1[5] ),
    .QN(_2991_));
 DFF_X1 \section_1.xn1[6]$_SDFF_PP0_  (.D(_0061_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\section_1.xn1[6] ),
    .QN(_2990_));
 DFF_X1 \section_1.xn1[7]$_SDFF_PP0_  (.D(_0062_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\section_1.xn1[7] ),
    .QN(_2989_));
 DFF_X1 \section_1.xn1[8]$_SDFF_PP0_  (.D(_0063_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\section_1.xn1[8] ),
    .QN(_2988_));
 DFF_X1 \section_1.xn1[9]$_SDFF_PP0_  (.D(_0064_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\section_1.xn1[9] ),
    .QN(_2987_));
 DFF_X1 \section_1.xn2[0]$_SDFF_PP0_  (.D(net13),
    .CK(clknet_3_1__leaf_clk),
    .Q(\section_1.xn2[0] ),
    .QN(_2986_));
 DFF_X1 \section_1.xn2[10]$_SDFF_PP0_  (.D(_0066_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\section_1.xn2[10] ),
    .QN(_2985_));
 DFF_X1 \section_1.xn2[1]$_SDFF_PP0_  (.D(net11),
    .CK(clknet_3_0__leaf_clk),
    .Q(\section_1.xn2[1] ),
    .QN(_2984_));
 DFF_X1 \section_1.xn2[2]$_SDFF_PP0_  (.D(net9),
    .CK(clknet_3_0__leaf_clk),
    .Q(\section_1.xn2[2] ),
    .QN(_2983_));
 DFF_X1 \section_1.xn2[3]$_SDFF_PP0_  (.D(net26),
    .CK(clknet_3_0__leaf_clk),
    .Q(\section_1.xn2[3] ),
    .QN(_2982_));
 DFF_X1 \section_1.xn2[4]$_SDFF_PP0_  (.D(_0070_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\section_1.xn2[4] ),
    .QN(_2981_));
 DFF_X1 \section_1.xn2[5]$_SDFF_PP0_  (.D(_0071_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\section_1.xn2[5] ),
    .QN(_2980_));
 DFF_X1 \section_1.xn2[6]$_SDFF_PP0_  (.D(net24),
    .CK(clknet_3_2__leaf_clk),
    .Q(\section_1.xn2[6] ),
    .QN(_2979_));
 DFF_X1 \section_1.xn2[7]$_SDFF_PP0_  (.D(net6),
    .CK(clknet_3_2__leaf_clk),
    .Q(\section_1.xn2[7] ),
    .QN(_2978_));
 DFF_X1 \section_1.xn2[8]$_SDFF_PP0_  (.D(net3),
    .CK(clknet_3_2__leaf_clk),
    .Q(\section_1.xn2[8] ),
    .QN(_2977_));
 DFF_X1 \section_1.xn2[9]$_SDFF_PP0_  (.D(_0075_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\section_1.xn2[9] ),
    .QN(_2976_));
 DFF_X1 \section_1.yn2[0]$_SDFF_PP0_  (.D(_0076_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\section_1.yn2[0] ),
    .QN(_0015_));
 DFF_X1 \section_1.yn2[10]$_SDFF_PP0_  (.D(_0077_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\section_1.yn2[10] ),
    .QN(_0004_));
 DFF_X1 \section_1.yn2[1]$_SDFF_PP0_  (.D(_0078_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\section_1.yn2[1] ),
    .QN(_0014_));
 DFF_X1 \section_1.yn2[2]$_SDFF_PP0_  (.D(_0079_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\section_1.yn2[2] ),
    .QN(_0013_));
 DFF_X1 \section_1.yn2[3]$_SDFF_PP0_  (.D(_0080_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\section_1.yn2[3] ),
    .QN(_0012_));
 DFF_X1 \section_1.yn2[4]$_SDFF_PP0_  (.D(_0081_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\section_1.yn2[4] ),
    .QN(_0011_));
 DFF_X1 \section_1.yn2[5]$_SDFF_PP0_  (.D(_0082_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\section_1.yn2[5] ),
    .QN(_0009_));
 DFF_X1 \section_1.yn2[6]$_SDFF_PP0_  (.D(_0083_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\section_1.yn2[6] ),
    .QN(_0003_));
 DFF_X1 \section_1.yn2[7]$_SDFF_PP0_  (.D(_0084_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\section_1.yn2[7] ),
    .QN(_0001_));
 DFF_X1 \section_1.yn2[8]$_SDFF_PP0_  (.D(_0085_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\section_1.yn2[8] ),
    .QN(_0008_));
 DFF_X1 \section_1.yn2[9]$_SDFF_PP0_  (.D(net68),
    .CK(clknet_3_3__leaf_clk),
    .Q(\section_1.yn2[9] ),
    .QN(_0030_));
 DFF_X1 \section_2.xn2[0]$_SDFF_PP0_  (.D(_0087_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\section_2.xn2[0] ),
    .QN(_0024_));
 DFF_X1 \section_2.xn2[10]$_SDFF_PP0_  (.D(_0088_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\section_2.xn2[10] ),
    .QN(_0031_));
 DFF_X1 \section_2.xn2[1]$_SDFF_PP0_  (.D(_0089_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\section_2.xn2[1] ),
    .QN(_0023_));
 DFF_X1 \section_2.xn2[2]$_SDFF_PP0_  (.D(_0090_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\section_2.xn2[2] ),
    .QN(_0022_));
 DFF_X1 \section_2.xn2[3]$_SDFF_PP0_  (.D(_0091_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\section_2.xn2[3] ),
    .QN(_0021_));
 DFF_X1 \section_2.xn2[4]$_SDFF_PP0_  (.D(_0092_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\section_2.xn2[4] ),
    .QN(_0019_));
 DFF_X1 \section_2.xn2[5]$_SDFF_PP0_  (.D(_0093_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\section_2.xn2[5] ),
    .QN(_0017_));
 DFF_X1 \section_2.xn2[6]$_SDFF_PP0_  (.D(_0094_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\section_2.xn2[6] ),
    .QN(_0020_));
 DFF_X1 \section_2.xn2[7]$_SDFF_PP0_  (.D(_0095_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\section_2.xn2[7] ),
    .QN(_0018_));
 DFF_X1 \section_2.xn2[8]$_SDFF_PP0_  (.D(_0096_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\section_2.xn2[8] ),
    .QN(_0016_));
 DFF_X1 \section_2.xn2[9]$_SDFF_PP0_  (.D(_0097_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\section_2.xn2[9] ),
    .QN(_2975_));
 DFF_X1 \section_2.yn2[0]$_SDFF_PP0_  (.D(_0098_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\section_2.yn2[0] ),
    .QN(_0029_));
 DFF_X1 \section_2.yn2[10]$_SDFF_PP0_  (.D(_0099_),
    .CK(clknet_3_7__leaf_clk),
    .Q(\section_2.yn2[10] ),
    .QN(_0002_));
 DFF_X1 \section_2.yn2[1]$_SDFF_PP0_  (.D(net55),
    .CK(clknet_3_5__leaf_clk),
    .Q(\section_2.yn2[1] ),
    .QN(_0027_));
 DFF_X1 \section_2.yn2[2]$_SDFF_PP0_  (.D(net57),
    .CK(clknet_3_5__leaf_clk),
    .Q(\section_2.yn2[2] ),
    .QN(_0025_));
 DFF_X1 \section_2.yn2[3]$_SDFF_PP0_  (.D(net51),
    .CK(clknet_3_5__leaf_clk),
    .Q(\section_2.yn2[3] ),
    .QN(_2974_));
 DFF_X1 \section_2.yn2[4]$_SDFF_PP0_  (.D(net53),
    .CK(clknet_3_5__leaf_clk),
    .Q(\section_2.yn2[4] ),
    .QN(_2973_));
 DFF_X1 \section_2.yn2[5]$_SDFF_PP0_  (.D(net49),
    .CK(clknet_3_5__leaf_clk),
    .Q(\section_2.yn2[5] ),
    .QN(_0028_));
 DFF_X1 \section_2.yn2[6]$_SDFF_PP0_  (.D(net76),
    .CK(clknet_3_7__leaf_clk),
    .Q(\section_2.yn2[6] ),
    .QN(_0026_));
 DFF_X1 \section_2.yn2[7]$_SDFF_PP0_  (.D(net59),
    .CK(clknet_3_7__leaf_clk),
    .Q(\section_2.yn2[7] ),
    .QN(_2972_));
 DFF_X1 \section_2.yn2[8]$_SDFF_PP0_  (.D(_0107_),
    .CK(clknet_3_7__leaf_clk),
    .Q(\section_2.yn2[8] ),
    .QN(_2971_));
 DFF_X1 \section_2.yn2[9]$_SDFF_PP0_  (.D(_0108_),
    .CK(clknet_3_7__leaf_clk),
    .Q(\section_2.yn2[9] ),
    .QN(_2970_));
 DFF_X1 \z[0]$_SDFF_PP0_  (.D(_0109_),
    .CK(clknet_3_5__leaf_clk),
    .Q(z[0]),
    .QN(_2969_));
 DFF_X1 \z[10]$_SDFF_PP0_  (.D(_0110_),
    .CK(clknet_3_7__leaf_clk),
    .Q(z[10]),
    .QN(_2968_));
 DFF_X1 \z[1]$_SDFF_PP0_  (.D(_0111_),
    .CK(clknet_3_5__leaf_clk),
    .Q(z[1]),
    .QN(_2967_));
 DFF_X1 \z[2]$_SDFF_PP0_  (.D(_0112_),
    .CK(clknet_3_5__leaf_clk),
    .Q(z[2]),
    .QN(_2966_));
 DFF_X1 \z[3]$_SDFF_PP0_  (.D(_0113_),
    .CK(clknet_3_5__leaf_clk),
    .Q(z[3]),
    .QN(_2965_));
 DFF_X1 \z[4]$_SDFF_PP0_  (.D(_0114_),
    .CK(clknet_3_5__leaf_clk),
    .Q(z[4]),
    .QN(_2964_));
 DFF_X1 \z[5]$_SDFF_PP0_  (.D(_0115_),
    .CK(clknet_3_7__leaf_clk),
    .Q(z[5]),
    .QN(_2963_));
 DFF_X1 \z[6]$_SDFF_PP0_  (.D(_0116_),
    .CK(clknet_3_7__leaf_clk),
    .Q(z[6]),
    .QN(_2962_));
 DFF_X1 \z[7]$_SDFF_PP0_  (.D(_0117_),
    .CK(clknet_3_7__leaf_clk),
    .Q(z[7]),
    .QN(_2961_));
 DFF_X1 \z[8]$_SDFF_PP0_  (.D(_0118_),
    .CK(clknet_3_7__leaf_clk),
    .Q(z[8]),
    .QN(_2960_));
 DFF_X1 \z[9]$_SDFF_PP0_  (.D(_0119_),
    .CK(clknet_3_7__leaf_clk),
    .Q(z[9]),
    .QN(_2959_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_103 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_104 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_105 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_106 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_107 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_108 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_109 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_110 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_111 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_112 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_113 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_114 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_115 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_116 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_117 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_118 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_119 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_120 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_121 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_122 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_123 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_124 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_125 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_126 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_127 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_128 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_129 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_130 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_131 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_132 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_133 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_134 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_135 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_136 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_137 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_138 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_139 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_140 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_141 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_142 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_143 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_144 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_145 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_146 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_147 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_148 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_149 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_150 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_151 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_152 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_153 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_154 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_155 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_156 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_157 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_158 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_159 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_160 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_161 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_162 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_163 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_164 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_165 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_166 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_167 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_168 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_169 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_170 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_171 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_172 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_173 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_174 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_175 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_176 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_177 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_178 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_179 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_180 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_181 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_182 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_183 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_184 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_185 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_186 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_187 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_41_188 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_41_189 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_190 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_191 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_43_192 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_43_193 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_194 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_195 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_45_196 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_45_197 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_198 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_199 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_47_200 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_47_201 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_202 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_203 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_49_204 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_49_205 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_206 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_207 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_208 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_209 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_210 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_211 ();
 CLKBUF_X1 hold1 (.A(\section_1.xn1[8] ),
    .Z(net1));
 CLKBUF_X1 hold2 (.A(_0921_),
    .Z(net2));
 CLKBUF_X1 hold3 (.A(_0074_),
    .Z(net3));
 CLKBUF_X1 hold4 (.A(\section_1.xn1[7] ),
    .Z(net4));
 CLKBUF_X1 hold5 (.A(_0922_),
    .Z(net5));
 CLKBUF_X1 hold6 (.A(_0073_),
    .Z(net6));
 CLKBUF_X1 hold7 (.A(\section_1.t1[2] ),
    .Z(net7));
 CLKBUF_X1 hold8 (.A(_0926_),
    .Z(net8));
 CLKBUF_X1 hold9 (.A(_0068_),
    .Z(net9));
 CLKBUF_X1 hold10 (.A(net94),
    .Z(net10));
 CLKBUF_X1 hold11 (.A(_0067_),
    .Z(net11));
 CLKBUF_X1 hold12 (.A(net93),
    .Z(net12));
 CLKBUF_X1 hold13 (.A(_0065_),
    .Z(net13));
 CLKBUF_X1 hold14 (.A(\in_reg1[10] ),
    .Z(net14));
 CLKBUF_X1 hold15 (.A(_0933_),
    .Z(net15));
 CLKBUF_X1 hold16 (.A(_0059_),
    .Z(net16));
 CLKBUF_X1 hold17 (.A(\in_reg1[5] ),
    .Z(net17));
 CLKBUF_X1 hold18 (.A(_0932_),
    .Z(net18));
 CLKBUF_X1 hold19 (.A(_0060_),
    .Z(net19));
 CLKBUF_X1 hold20 (.A(net104),
    .Z(net20));
 CLKBUF_X1 hold21 (.A(_0920_),
    .Z(net21));
 CLKBUF_X1 hold22 (.A(\section_1.xn1[6] ),
    .Z(net22));
 CLKBUF_X1 hold23 (.A(_0923_),
    .Z(net23));
 CLKBUF_X1 hold24 (.A(_0072_),
    .Z(net24));
 CLKBUF_X1 hold25 (.A(net95),
    .Z(net25));
 CLKBUF_X1 hold26 (.A(_0069_),
    .Z(net26));
 CLKBUF_X1 hold27 (.A(net100),
    .Z(net27));
 CLKBUF_X1 hold28 (.A(_0925_),
    .Z(net28));
 CLKBUF_X1 hold29 (.A(net96),
    .Z(net29));
 CLKBUF_X1 hold30 (.A(_0054_),
    .Z(net30));
 CLKBUF_X1 hold31 (.A(net105),
    .Z(net31));
 CLKBUF_X1 hold32 (.A(_0934_),
    .Z(net32));
 CLKBUF_X1 hold33 (.A(net110),
    .Z(net33));
 CLKBUF_X1 hold34 (.A(_0928_),
    .Z(net34));
 CLKBUF_X1 hold35 (.A(net111),
    .Z(net35));
 CLKBUF_X1 hold36 (.A(_0929_),
    .Z(net36));
 CLKBUF_X1 hold37 (.A(net108),
    .Z(net37));
 CLKBUF_X1 hold38 (.A(_0931_),
    .Z(net38));
 CLKBUF_X1 hold39 (.A(net109),
    .Z(net39));
 CLKBUF_X1 hold40 (.A(_0924_),
    .Z(net40));
 CLKBUF_X1 hold41 (.A(net115),
    .Z(net41));
 CLKBUF_X1 hold42 (.A(_2386_),
    .Z(net42));
 CLKBUF_X1 hold43 (.A(net122),
    .Z(net43));
 CLKBUF_X1 hold44 (.A(_0930_),
    .Z(net44));
 CLKBUF_X1 hold45 (.A(\in_reg1[2] ),
    .Z(net45));
 CLKBUF_X1 hold46 (.A(_0936_),
    .Z(net46));
 CLKBUF_X1 hold47 (.A(net97),
    .Z(net47));
 CLKBUF_X1 hold48 (.A(net114),
    .Z(net48));
 CLKBUF_X1 hold49 (.A(_0104_),
    .Z(net49));
 CLKBUF_X1 hold50 (.A(net118),
    .Z(net50));
 CLKBUF_X1 hold51 (.A(_0102_),
    .Z(net51));
 CLKBUF_X1 hold52 (.A(net121),
    .Z(net52));
 CLKBUF_X1 hold53 (.A(_0103_),
    .Z(net53));
 CLKBUF_X1 hold54 (.A(net120),
    .Z(net54));
 CLKBUF_X1 hold55 (.A(_0100_),
    .Z(net55));
 CLKBUF_X1 hold56 (.A(net119),
    .Z(net56));
 CLKBUF_X1 hold57 (.A(_0101_),
    .Z(net57));
 CLKBUF_X1 hold58 (.A(net123),
    .Z(net58));
 CLKBUF_X1 hold59 (.A(_0106_),
    .Z(net59));
 CLKBUF_X1 hold60 (.A(z[0]),
    .Z(net60));
 CLKBUF_X1 hold61 (.A(_2862_),
    .Z(net61));
 CLKBUF_X1 hold62 (.A(net98),
    .Z(net62));
 CLKBUF_X1 hold63 (.A(\section_1.yn2[6] ),
    .Z(net63));
 CLKBUF_X1 hold64 (.A(_2328_),
    .Z(net64));
 CLKBUF_X1 hold65 (.A(\section_1.yn2[3] ),
    .Z(net65));
 CLKBUF_X1 hold66 (.A(_0917_),
    .Z(net66));
 CLKBUF_X1 hold67 (.A(\coll_reg[9] ),
    .Z(net67));
 CLKBUF_X1 hold68 (.A(_0086_),
    .Z(net68));
 CLKBUF_X1 hold69 (.A(z[9]),
    .Z(net69));
 CLKBUF_X1 hold70 (.A(_2767_),
    .Z(net70));
 CLKBUF_X1 hold71 (.A(\section_1.yn2[2] ),
    .Z(net71));
 CLKBUF_X1 hold72 (.A(_1528_),
    .Z(net72));
 CLKBUF_X1 hold73 (.A(\section_1.xn1[10] ),
    .Z(net73));
 CLKBUF_X1 hold74 (.A(_0927_),
    .Z(net74));
 CLKBUF_X1 hold75 (.A(z[6]),
    .Z(net75));
 CLKBUF_X1 hold76 (.A(_0105_),
    .Z(net76));
 CLKBUF_X1 hold77 (.A(\section_1.yn2[8] ),
    .Z(net77));
 CLKBUF_X1 hold78 (.A(_2504_),
    .Z(net78));
 CLKBUF_X1 hold79 (.A(net101),
    .Z(net79));
 CLKBUF_X1 hold80 (.A(net99),
    .Z(net80));
 CLKBUF_X1 hold81 (.A(net102),
    .Z(net81));
 CLKBUF_X1 hold82 (.A(net103),
    .Z(net82));
 CLKBUF_X1 hold83 (.A(net106),
    .Z(net83));
 CLKBUF_X1 hold84 (.A(net107),
    .Z(net84));
 CLKBUF_X1 hold85 (.A(net112),
    .Z(net85));
 CLKBUF_X1 hold86 (.A(net117),
    .Z(net86));
 CLKBUF_X1 hold87 (.A(\coll_reg[5] ),
    .Z(net87));
 CLKBUF_X1 hold88 (.A(\coll_reg[6] ),
    .Z(net88));
 CLKBUF_X1 hold89 (.A(\coll_reg[10] ),
    .Z(net89));
 CLKBUF_X1 hold90 (.A(\coll_reg[4] ),
    .Z(net90));
 CLKBUF_X1 hold91 (.A(\coll_reg[3] ),
    .Z(net91));
 CLKBUF_X1 hold92 (.A(\coll_reg[8] ),
    .Z(net92));
 CLKBUF_X1 hold93 (.A(\section_1.t1[0] ),
    .Z(net93));
 CLKBUF_X1 hold94 (.A(\section_1.t1[1] ),
    .Z(net94));
 CLKBUF_X1 hold95 (.A(\section_1.t1[3] ),
    .Z(net95));
 CLKBUF_X1 hold96 (.A(\in_reg1[0] ),
    .Z(net96));
 BUF_X8 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 BUF_X8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_0__leaf_clk));
 BUF_X8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_1__leaf_clk));
 BUF_X8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_2__leaf_clk));
 BUF_X8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_3__leaf_clk));
 BUF_X8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_4__leaf_clk));
 BUF_X8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_5__leaf_clk));
 BUF_X8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_6__leaf_clk));
 BUF_X8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_7__leaf_clk));
 BUF_X8 clkload0 (.A(clknet_3_1__leaf_clk));
 INV_X2 clkload1 (.A(clknet_3_2__leaf_clk));
 BUF_X8 clkload2 (.A(clknet_3_3__leaf_clk));
 BUF_X8 clkload3 (.A(clknet_3_4__leaf_clk));
 BUF_X4 clkload4 (.A(clknet_3_5__leaf_clk));
 BUF_X8 clkload5 (.A(clknet_3_6__leaf_clk));
 BUF_X4 clkload6 (.A(clknet_3_7__leaf_clk));
 CLKBUF_X1 hold97 (.A(\in_reg1[3] ),
    .Z(net97));
 CLKBUF_X1 hold98 (.A(\in_reg1[1] ),
    .Z(net98));
 CLKBUF_X1 hold99 (.A(\section_1.yn2[4] ),
    .Z(net99));
 CLKBUF_X1 hold100 (.A(\section_1.t1[4] ),
    .Z(net100));
 CLKBUF_X1 hold101 (.A(z[8]),
    .Z(net101));
 CLKBUF_X1 hold102 (.A(z[10]),
    .Z(net102));
 CLKBUF_X1 hold103 (.A(\section_1.yn2[1] ),
    .Z(net103));
 CLKBUF_X1 hold104 (.A(\section_1.xn1[9] ),
    .Z(net104));
 CLKBUF_X1 hold105 (.A(\in_reg1[4] ),
    .Z(net105));
 CLKBUF_X1 hold106 (.A(\section_1.yn2[9] ),
    .Z(net106));
 CLKBUF_X1 hold107 (.A(\coll_reg[2] ),
    .Z(net107));
 CLKBUF_X1 hold108 (.A(\in_reg1[6] ),
    .Z(net108));
 CLKBUF_X1 hold109 (.A(\section_1.xn1[5] ),
    .Z(net109));
 CLKBUF_X1 hold110 (.A(\in_reg1[9] ),
    .Z(net110));
 CLKBUF_X1 hold111 (.A(\in_reg1[8] ),
    .Z(net111));
 CLKBUF_X1 hold112 (.A(\section_1.yn2[7] ),
    .Z(net112));
 CLKBUF_X1 hold113 (.A(\coll_reg[7] ),
    .Z(net113));
 CLKBUF_X1 hold114 (.A(z[5]),
    .Z(net114));
 CLKBUF_X1 hold115 (.A(\section_1.yn2[0] ),
    .Z(net115));
 CLKBUF_X1 hold116 (.A(\coll_reg[1] ),
    .Z(net116));
 CLKBUF_X1 hold117 (.A(\section_1.yn2[5] ),
    .Z(net117));
 CLKBUF_X1 hold118 (.A(z[3]),
    .Z(net118));
 CLKBUF_X1 hold119 (.A(z[2]),
    .Z(net119));
 CLKBUF_X1 hold120 (.A(z[1]),
    .Z(net120));
 CLKBUF_X1 hold121 (.A(z[4]),
    .Z(net121));
 CLKBUF_X1 hold122 (.A(\in_reg1[7] ),
    .Z(net122));
 CLKBUF_X1 hold123 (.A(z[7]),
    .Z(net123));
 FILLCELL_X16 FILLER_0_0_1 ();
 FILLCELL_X2 FILLER_0_0_17 ();
 FILLCELL_X1 FILLER_0_0_19 ();
 FILLCELL_X8 FILLER_0_0_22 ();
 FILLCELL_X4 FILLER_0_0_34 ();
 FILLCELL_X2 FILLER_0_0_75 ();
 FILLCELL_X8 FILLER_0_0_81 ();
 FILLCELL_X4 FILLER_0_0_90 ();
 FILLCELL_X2 FILLER_0_0_94 ();
 FILLCELL_X1 FILLER_0_0_96 ();
 FILLCELL_X2 FILLER_0_0_100 ();
 FILLCELL_X1 FILLER_0_0_102 ();
 FILLCELL_X4 FILLER_0_0_106 ();
 FILLCELL_X1 FILLER_0_0_110 ();
 FILLCELL_X4 FILLER_0_0_131 ();
 FILLCELL_X1 FILLER_0_0_135 ();
 FILLCELL_X1 FILLER_0_0_153 ();
 FILLCELL_X1 FILLER_0_0_157 ();
 FILLCELL_X1 FILLER_0_0_162 ();
 FILLCELL_X1 FILLER_0_0_167 ();
 FILLCELL_X1 FILLER_0_0_171 ();
 FILLCELL_X1 FILLER_0_0_177 ();
 FILLCELL_X2 FILLER_0_0_181 ();
 FILLCELL_X1 FILLER_0_0_186 ();
 FILLCELL_X1 FILLER_0_0_191 ();
 FILLCELL_X2 FILLER_0_0_197 ();
 FILLCELL_X8 FILLER_0_0_203 ();
 FILLCELL_X4 FILLER_0_0_211 ();
 FILLCELL_X1 FILLER_0_0_215 ();
 FILLCELL_X1 FILLER_0_0_240 ();
 FILLCELL_X1 FILLER_0_0_257 ();
 FILLCELL_X2 FILLER_0_0_271 ();
 FILLCELL_X16 FILLER_0_0_293 ();
 FILLCELL_X4 FILLER_0_0_309 ();
 FILLCELL_X8 FILLER_0_0_319 ();
 FILLCELL_X4 FILLER_0_0_327 ();
 FILLCELL_X4 FILLER_0_0_334 ();
 FILLCELL_X4 FILLER_0_0_344 ();
 FILLCELL_X2 FILLER_0_0_348 ();
 FILLCELL_X1 FILLER_0_0_357 ();
 FILLCELL_X16 FILLER_0_0_361 ();
 FILLCELL_X8 FILLER_0_0_377 ();
 FILLCELL_X2 FILLER_0_0_385 ();
 FILLCELL_X1 FILLER_0_0_387 ();
 FILLCELL_X32 FILLER_0_1_1 ();
 FILLCELL_X8 FILLER_0_1_33 ();
 FILLCELL_X2 FILLER_0_1_41 ();
 FILLCELL_X2 FILLER_0_1_46 ();
 FILLCELL_X1 FILLER_0_1_48 ();
 FILLCELL_X2 FILLER_0_1_52 ();
 FILLCELL_X1 FILLER_0_1_54 ();
 FILLCELL_X1 FILLER_0_1_149 ();
 FILLCELL_X1 FILLER_0_1_212 ();
 FILLCELL_X1 FILLER_0_1_223 ();
 FILLCELL_X1 FILLER_0_1_258 ();
 FILLCELL_X1 FILLER_0_1_276 ();
 FILLCELL_X1 FILLER_0_1_279 ();
 FILLCELL_X1 FILLER_0_1_331 ();
 FILLCELL_X2 FILLER_0_1_348 ();
 FILLCELL_X1 FILLER_0_1_352 ();
 FILLCELL_X8 FILLER_0_1_378 ();
 FILLCELL_X2 FILLER_0_1_386 ();
 FILLCELL_X32 FILLER_0_2_1 ();
 FILLCELL_X1 FILLER_0_2_33 ();
 FILLCELL_X1 FILLER_0_2_37 ();
 FILLCELL_X2 FILLER_0_2_67 ();
 FILLCELL_X2 FILLER_0_2_94 ();
 FILLCELL_X2 FILLER_0_2_102 ();
 FILLCELL_X1 FILLER_0_2_129 ();
 FILLCELL_X1 FILLER_0_2_133 ();
 FILLCELL_X2 FILLER_0_2_149 ();
 FILLCELL_X1 FILLER_0_2_160 ();
 FILLCELL_X1 FILLER_0_2_164 ();
 FILLCELL_X1 FILLER_0_2_171 ();
 FILLCELL_X1 FILLER_0_2_176 ();
 FILLCELL_X1 FILLER_0_2_180 ();
 FILLCELL_X1 FILLER_0_2_187 ();
 FILLCELL_X1 FILLER_0_2_192 ();
 FILLCELL_X1 FILLER_0_2_245 ();
 FILLCELL_X1 FILLER_0_2_260 ();
 FILLCELL_X4 FILLER_0_2_268 ();
 FILLCELL_X1 FILLER_0_2_272 ();
 FILLCELL_X2 FILLER_0_2_287 ();
 FILLCELL_X1 FILLER_0_2_289 ();
 FILLCELL_X1 FILLER_0_2_293 ();
 FILLCELL_X1 FILLER_0_2_298 ();
 FILLCELL_X1 FILLER_0_2_316 ();
 FILLCELL_X2 FILLER_0_2_360 ();
 FILLCELL_X1 FILLER_0_2_377 ();
 FILLCELL_X4 FILLER_0_2_383 ();
 FILLCELL_X1 FILLER_0_2_387 ();
 FILLCELL_X16 FILLER_0_3_1 ();
 FILLCELL_X2 FILLER_0_3_17 ();
 FILLCELL_X8 FILLER_0_3_39 ();
 FILLCELL_X2 FILLER_0_3_47 ();
 FILLCELL_X2 FILLER_0_3_79 ();
 FILLCELL_X4 FILLER_0_3_94 ();
 FILLCELL_X2 FILLER_0_3_98 ();
 FILLCELL_X1 FILLER_0_3_100 ();
 FILLCELL_X1 FILLER_0_3_140 ();
 FILLCELL_X2 FILLER_0_3_144 ();
 FILLCELL_X1 FILLER_0_3_158 ();
 FILLCELL_X1 FILLER_0_3_162 ();
 FILLCELL_X1 FILLER_0_3_166 ();
 FILLCELL_X2 FILLER_0_3_170 ();
 FILLCELL_X4 FILLER_0_3_189 ();
 FILLCELL_X2 FILLER_0_3_193 ();
 FILLCELL_X1 FILLER_0_3_195 ();
 FILLCELL_X1 FILLER_0_3_202 ();
 FILLCELL_X1 FILLER_0_3_218 ();
 FILLCELL_X1 FILLER_0_3_222 ();
 FILLCELL_X2 FILLER_0_3_225 ();
 FILLCELL_X1 FILLER_0_3_232 ();
 FILLCELL_X2 FILLER_0_3_236 ();
 FILLCELL_X2 FILLER_0_3_241 ();
 FILLCELL_X1 FILLER_0_3_243 ();
 FILLCELL_X1 FILLER_0_3_250 ();
 FILLCELL_X2 FILLER_0_3_267 ();
 FILLCELL_X4 FILLER_0_3_289 ();
 FILLCELL_X1 FILLER_0_3_293 ();
 FILLCELL_X1 FILLER_0_3_307 ();
 FILLCELL_X2 FILLER_0_3_317 ();
 FILLCELL_X1 FILLER_0_3_365 ();
 FILLCELL_X1 FILLER_0_3_370 ();
 FILLCELL_X8 FILLER_0_3_376 ();
 FILLCELL_X4 FILLER_0_3_384 ();
 FILLCELL_X16 FILLER_0_4_1 ();
 FILLCELL_X8 FILLER_0_4_17 ();
 FILLCELL_X2 FILLER_0_4_35 ();
 FILLCELL_X4 FILLER_0_4_60 ();
 FILLCELL_X1 FILLER_0_4_64 ();
 FILLCELL_X2 FILLER_0_4_81 ();
 FILLCELL_X2 FILLER_0_4_99 ();
 FILLCELL_X4 FILLER_0_4_104 ();
 FILLCELL_X2 FILLER_0_4_131 ();
 FILLCELL_X1 FILLER_0_4_135 ();
 FILLCELL_X2 FILLER_0_4_146 ();
 FILLCELL_X2 FILLER_0_4_151 ();
 FILLCELL_X2 FILLER_0_4_157 ();
 FILLCELL_X2 FILLER_0_4_163 ();
 FILLCELL_X1 FILLER_0_4_165 ();
 FILLCELL_X2 FILLER_0_4_169 ();
 FILLCELL_X1 FILLER_0_4_171 ();
 FILLCELL_X2 FILLER_0_4_178 ();
 FILLCELL_X8 FILLER_0_4_203 ();
 FILLCELL_X2 FILLER_0_4_211 ();
 FILLCELL_X1 FILLER_0_4_213 ();
 FILLCELL_X1 FILLER_0_4_287 ();
 FILLCELL_X4 FILLER_0_4_297 ();
 FILLCELL_X2 FILLER_0_4_301 ();
 FILLCELL_X1 FILLER_0_4_303 ();
 FILLCELL_X2 FILLER_0_4_323 ();
 FILLCELL_X1 FILLER_0_4_325 ();
 FILLCELL_X1 FILLER_0_4_334 ();
 FILLCELL_X1 FILLER_0_4_339 ();
 FILLCELL_X1 FILLER_0_4_343 ();
 FILLCELL_X4 FILLER_0_4_350 ();
 FILLCELL_X2 FILLER_0_4_354 ();
 FILLCELL_X8 FILLER_0_4_360 ();
 FILLCELL_X1 FILLER_0_4_368 ();
 FILLCELL_X2 FILLER_0_4_386 ();
 FILLCELL_X4 FILLER_0_5_1 ();
 FILLCELL_X2 FILLER_0_5_39 ();
 FILLCELL_X4 FILLER_0_5_53 ();
 FILLCELL_X1 FILLER_0_5_72 ();
 FILLCELL_X1 FILLER_0_5_76 ();
 FILLCELL_X1 FILLER_0_5_87 ();
 FILLCELL_X1 FILLER_0_5_91 ();
 FILLCELL_X1 FILLER_0_5_98 ();
 FILLCELL_X1 FILLER_0_5_103 ();
 FILLCELL_X1 FILLER_0_5_110 ();
 FILLCELL_X2 FILLER_0_5_130 ();
 FILLCELL_X1 FILLER_0_5_135 ();
 FILLCELL_X2 FILLER_0_5_156 ();
 FILLCELL_X1 FILLER_0_5_170 ();
 FILLCELL_X2 FILLER_0_5_175 ();
 FILLCELL_X1 FILLER_0_5_177 ();
 FILLCELL_X4 FILLER_0_5_199 ();
 FILLCELL_X1 FILLER_0_5_209 ();
 FILLCELL_X1 FILLER_0_5_213 ();
 FILLCELL_X2 FILLER_0_5_220 ();
 FILLCELL_X2 FILLER_0_5_225 ();
 FILLCELL_X8 FILLER_0_5_230 ();
 FILLCELL_X2 FILLER_0_5_240 ();
 FILLCELL_X1 FILLER_0_5_244 ();
 FILLCELL_X2 FILLER_0_5_251 ();
 FILLCELL_X1 FILLER_0_5_271 ();
 FILLCELL_X2 FILLER_0_5_276 ();
 FILLCELL_X2 FILLER_0_5_293 ();
 FILLCELL_X1 FILLER_0_5_304 ();
 FILLCELL_X1 FILLER_0_5_309 ();
 FILLCELL_X2 FILLER_0_5_317 ();
 FILLCELL_X1 FILLER_0_5_328 ();
 FILLCELL_X1 FILLER_0_5_370 ();
 FILLCELL_X4 FILLER_0_6_1 ();
 FILLCELL_X2 FILLER_0_6_5 ();
 FILLCELL_X8 FILLER_0_6_11 ();
 FILLCELL_X2 FILLER_0_6_19 ();
 FILLCELL_X2 FILLER_0_6_25 ();
 FILLCELL_X2 FILLER_0_6_49 ();
 FILLCELL_X4 FILLER_0_6_60 ();
 FILLCELL_X1 FILLER_0_6_64 ();
 FILLCELL_X4 FILLER_0_6_84 ();
 FILLCELL_X1 FILLER_0_6_88 ();
 FILLCELL_X1 FILLER_0_6_90 ();
 FILLCELL_X1 FILLER_0_6_109 ();
 FILLCELL_X4 FILLER_0_6_115 ();
 FILLCELL_X1 FILLER_0_6_119 ();
 FILLCELL_X2 FILLER_0_6_138 ();
 FILLCELL_X2 FILLER_0_6_159 ();
 FILLCELL_X1 FILLER_0_6_170 ();
 FILLCELL_X4 FILLER_0_6_174 ();
 FILLCELL_X2 FILLER_0_6_180 ();
 FILLCELL_X1 FILLER_0_6_182 ();
 FILLCELL_X4 FILLER_0_6_237 ();
 FILLCELL_X1 FILLER_0_6_241 ();
 FILLCELL_X4 FILLER_0_6_246 ();
 FILLCELL_X1 FILLER_0_6_250 ();
 FILLCELL_X2 FILLER_0_6_268 ();
 FILLCELL_X1 FILLER_0_6_284 ();
 FILLCELL_X8 FILLER_0_6_290 ();
 FILLCELL_X1 FILLER_0_6_298 ();
 FILLCELL_X1 FILLER_0_6_320 ();
 FILLCELL_X16 FILLER_0_6_328 ();
 FILLCELL_X4 FILLER_0_6_344 ();
 FILLCELL_X1 FILLER_0_6_369 ();
 FILLCELL_X8 FILLER_0_6_377 ();
 FILLCELL_X2 FILLER_0_6_385 ();
 FILLCELL_X1 FILLER_0_6_387 ();
 FILLCELL_X4 FILLER_0_7_1 ();
 FILLCELL_X2 FILLER_0_7_5 ();
 FILLCELL_X1 FILLER_0_7_24 ();
 FILLCELL_X1 FILLER_0_7_28 ();
 FILLCELL_X1 FILLER_0_7_39 ();
 FILLCELL_X1 FILLER_0_7_61 ();
 FILLCELL_X1 FILLER_0_7_68 ();
 FILLCELL_X1 FILLER_0_7_80 ();
 FILLCELL_X2 FILLER_0_7_102 ();
 FILLCELL_X2 FILLER_0_7_107 ();
 FILLCELL_X1 FILLER_0_7_113 ();
 FILLCELL_X4 FILLER_0_7_117 ();
 FILLCELL_X1 FILLER_0_7_134 ();
 FILLCELL_X2 FILLER_0_7_139 ();
 FILLCELL_X2 FILLER_0_7_147 ();
 FILLCELL_X2 FILLER_0_7_155 ();
 FILLCELL_X1 FILLER_0_7_157 ();
 FILLCELL_X1 FILLER_0_7_164 ();
 FILLCELL_X1 FILLER_0_7_169 ();
 FILLCELL_X1 FILLER_0_7_189 ();
 FILLCELL_X2 FILLER_0_7_196 ();
 FILLCELL_X1 FILLER_0_7_202 ();
 FILLCELL_X2 FILLER_0_7_209 ();
 FILLCELL_X4 FILLER_0_7_240 ();
 FILLCELL_X1 FILLER_0_7_244 ();
 FILLCELL_X2 FILLER_0_7_254 ();
 FILLCELL_X1 FILLER_0_7_256 ();
 FILLCELL_X1 FILLER_0_7_263 ();
 FILLCELL_X4 FILLER_0_7_270 ();
 FILLCELL_X1 FILLER_0_7_274 ();
 FILLCELL_X2 FILLER_0_7_280 ();
 FILLCELL_X1 FILLER_0_7_282 ();
 FILLCELL_X2 FILLER_0_7_287 ();
 FILLCELL_X2 FILLER_0_7_292 ();
 FILLCELL_X8 FILLER_0_7_306 ();
 FILLCELL_X4 FILLER_0_7_314 ();
 FILLCELL_X1 FILLER_0_7_318 ();
 FILLCELL_X8 FILLER_0_7_327 ();
 FILLCELL_X4 FILLER_0_7_335 ();
 FILLCELL_X4 FILLER_0_7_345 ();
 FILLCELL_X1 FILLER_0_7_349 ();
 FILLCELL_X1 FILLER_0_7_370 ();
 FILLCELL_X4 FILLER_0_8_1 ();
 FILLCELL_X1 FILLER_0_8_5 ();
 FILLCELL_X2 FILLER_0_8_41 ();
 FILLCELL_X2 FILLER_0_8_54 ();
 FILLCELL_X1 FILLER_0_8_69 ();
 FILLCELL_X1 FILLER_0_8_88 ();
 FILLCELL_X1 FILLER_0_8_90 ();
 FILLCELL_X2 FILLER_0_8_119 ();
 FILLCELL_X8 FILLER_0_8_131 ();
 FILLCELL_X4 FILLER_0_8_139 ();
 FILLCELL_X1 FILLER_0_8_143 ();
 FILLCELL_X2 FILLER_0_8_155 ();
 FILLCELL_X1 FILLER_0_8_166 ();
 FILLCELL_X4 FILLER_0_8_213 ();
 FILLCELL_X2 FILLER_0_8_217 ();
 FILLCELL_X16 FILLER_0_8_224 ();
 FILLCELL_X2 FILLER_0_8_240 ();
 FILLCELL_X2 FILLER_0_8_255 ();
 FILLCELL_X1 FILLER_0_8_260 ();
 FILLCELL_X8 FILLER_0_8_268 ();
 FILLCELL_X4 FILLER_0_8_276 ();
 FILLCELL_X1 FILLER_0_8_280 ();
 FILLCELL_X2 FILLER_0_8_287 ();
 FILLCELL_X2 FILLER_0_8_293 ();
 FILLCELL_X1 FILLER_0_8_295 ();
 FILLCELL_X1 FILLER_0_8_305 ();
 FILLCELL_X4 FILLER_0_8_315 ();
 FILLCELL_X1 FILLER_0_8_325 ();
 FILLCELL_X4 FILLER_0_8_329 ();
 FILLCELL_X1 FILLER_0_8_333 ();
 FILLCELL_X1 FILLER_0_8_353 ();
 FILLCELL_X2 FILLER_0_8_357 ();
 FILLCELL_X2 FILLER_0_8_365 ();
 FILLCELL_X2 FILLER_0_8_371 ();
 FILLCELL_X1 FILLER_0_8_373 ();
 FILLCELL_X8 FILLER_0_8_378 ();
 FILLCELL_X2 FILLER_0_8_386 ();
 FILLCELL_X4 FILLER_0_9_1 ();
 FILLCELL_X1 FILLER_0_9_14 ();
 FILLCELL_X1 FILLER_0_9_34 ();
 FILLCELL_X1 FILLER_0_9_37 ();
 FILLCELL_X4 FILLER_0_9_50 ();
 FILLCELL_X2 FILLER_0_9_57 ();
 FILLCELL_X1 FILLER_0_9_59 ();
 FILLCELL_X8 FILLER_0_9_69 ();
 FILLCELL_X1 FILLER_0_9_77 ();
 FILLCELL_X8 FILLER_0_9_91 ();
 FILLCELL_X4 FILLER_0_9_99 ();
 FILLCELL_X4 FILLER_0_9_118 ();
 FILLCELL_X1 FILLER_0_9_122 ();
 FILLCELL_X2 FILLER_0_9_135 ();
 FILLCELL_X1 FILLER_0_9_137 ();
 FILLCELL_X8 FILLER_0_9_153 ();
 FILLCELL_X4 FILLER_0_9_161 ();
 FILLCELL_X1 FILLER_0_9_165 ();
 FILLCELL_X4 FILLER_0_9_179 ();
 FILLCELL_X8 FILLER_0_9_187 ();
 FILLCELL_X4 FILLER_0_9_195 ();
 FILLCELL_X2 FILLER_0_9_199 ();
 FILLCELL_X1 FILLER_0_9_201 ();
 FILLCELL_X2 FILLER_0_9_218 ();
 FILLCELL_X4 FILLER_0_9_224 ();
 FILLCELL_X2 FILLER_0_9_238 ();
 FILLCELL_X1 FILLER_0_9_240 ();
 FILLCELL_X1 FILLER_0_9_247 ();
 FILLCELL_X1 FILLER_0_9_252 ();
 FILLCELL_X1 FILLER_0_9_262 ();
 FILLCELL_X2 FILLER_0_9_282 ();
 FILLCELL_X2 FILLER_0_9_310 ();
 FILLCELL_X2 FILLER_0_9_334 ();
 FILLCELL_X2 FILLER_0_9_360 ();
 FILLCELL_X16 FILLER_0_9_370 ();
 FILLCELL_X2 FILLER_0_9_386 ();
 FILLCELL_X8 FILLER_0_10_1 ();
 FILLCELL_X2 FILLER_0_10_9 ();
 FILLCELL_X2 FILLER_0_10_14 ();
 FILLCELL_X1 FILLER_0_10_16 ();
 FILLCELL_X2 FILLER_0_10_38 ();
 FILLCELL_X1 FILLER_0_10_50 ();
 FILLCELL_X1 FILLER_0_10_65 ();
 FILLCELL_X8 FILLER_0_10_74 ();
 FILLCELL_X2 FILLER_0_10_82 ();
 FILLCELL_X1 FILLER_0_10_84 ();
 FILLCELL_X16 FILLER_0_10_90 ();
 FILLCELL_X4 FILLER_0_10_106 ();
 FILLCELL_X1 FILLER_0_10_110 ();
 FILLCELL_X8 FILLER_0_10_115 ();
 FILLCELL_X1 FILLER_0_10_123 ();
 FILLCELL_X1 FILLER_0_10_130 ();
 FILLCELL_X1 FILLER_0_10_135 ();
 FILLCELL_X1 FILLER_0_10_142 ();
 FILLCELL_X2 FILLER_0_10_146 ();
 FILLCELL_X1 FILLER_0_10_194 ();
 FILLCELL_X2 FILLER_0_10_198 ();
 FILLCELL_X1 FILLER_0_10_213 ();
 FILLCELL_X1 FILLER_0_10_218 ();
 FILLCELL_X1 FILLER_0_10_223 ();
 FILLCELL_X2 FILLER_0_10_228 ();
 FILLCELL_X1 FILLER_0_10_240 ();
 FILLCELL_X1 FILLER_0_10_248 ();
 FILLCELL_X4 FILLER_0_10_259 ();
 FILLCELL_X4 FILLER_0_10_279 ();
 FILLCELL_X2 FILLER_0_10_283 ();
 FILLCELL_X8 FILLER_0_10_295 ();
 FILLCELL_X2 FILLER_0_10_312 ();
 FILLCELL_X1 FILLER_0_10_314 ();
 FILLCELL_X1 FILLER_0_10_321 ();
 FILLCELL_X1 FILLER_0_10_328 ();
 FILLCELL_X1 FILLER_0_10_332 ();
 FILLCELL_X1 FILLER_0_10_339 ();
 FILLCELL_X1 FILLER_0_10_343 ();
 FILLCELL_X1 FILLER_0_10_350 ();
 FILLCELL_X2 FILLER_0_10_356 ();
 FILLCELL_X2 FILLER_0_10_375 ();
 FILLCELL_X1 FILLER_0_10_387 ();
 FILLCELL_X4 FILLER_0_11_1 ();
 FILLCELL_X2 FILLER_0_11_5 ();
 FILLCELL_X1 FILLER_0_11_7 ();
 FILLCELL_X4 FILLER_0_11_34 ();
 FILLCELL_X1 FILLER_0_11_38 ();
 FILLCELL_X8 FILLER_0_11_42 ();
 FILLCELL_X4 FILLER_0_11_50 ();
 FILLCELL_X2 FILLER_0_11_60 ();
 FILLCELL_X2 FILLER_0_11_64 ();
 FILLCELL_X4 FILLER_0_11_76 ();
 FILLCELL_X2 FILLER_0_11_83 ();
 FILLCELL_X1 FILLER_0_11_91 ();
 FILLCELL_X1 FILLER_0_11_98 ();
 FILLCELL_X1 FILLER_0_11_102 ();
 FILLCELL_X1 FILLER_0_11_107 ();
 FILLCELL_X8 FILLER_0_11_149 ();
 FILLCELL_X8 FILLER_0_11_167 ();
 FILLCELL_X2 FILLER_0_11_175 ();
 FILLCELL_X1 FILLER_0_11_177 ();
 FILLCELL_X2 FILLER_0_11_182 ();
 FILLCELL_X1 FILLER_0_11_184 ();
 FILLCELL_X1 FILLER_0_11_189 ();
 FILLCELL_X1 FILLER_0_11_193 ();
 FILLCELL_X1 FILLER_0_11_197 ();
 FILLCELL_X2 FILLER_0_11_202 ();
 FILLCELL_X1 FILLER_0_11_253 ();
 FILLCELL_X1 FILLER_0_11_261 ();
 FILLCELL_X4 FILLER_0_11_265 ();
 FILLCELL_X2 FILLER_0_11_269 ();
 FILLCELL_X1 FILLER_0_11_280 ();
 FILLCELL_X1 FILLER_0_11_284 ();
 FILLCELL_X1 FILLER_0_11_294 ();
 FILLCELL_X8 FILLER_0_11_311 ();
 FILLCELL_X1 FILLER_0_11_319 ();
 FILLCELL_X2 FILLER_0_11_342 ();
 FILLCELL_X1 FILLER_0_11_344 ();
 FILLCELL_X1 FILLER_0_11_355 ();
 FILLCELL_X4 FILLER_0_11_363 ();
 FILLCELL_X1 FILLER_0_11_381 ();
 FILLCELL_X2 FILLER_0_11_385 ();
 FILLCELL_X1 FILLER_0_11_387 ();
 FILLCELL_X4 FILLER_0_12_1 ();
 FILLCELL_X2 FILLER_0_12_5 ();
 FILLCELL_X8 FILLER_0_12_11 ();
 FILLCELL_X2 FILLER_0_12_19 ();
 FILLCELL_X1 FILLER_0_12_21 ();
 FILLCELL_X1 FILLER_0_12_35 ();
 FILLCELL_X2 FILLER_0_12_56 ();
 FILLCELL_X2 FILLER_0_12_74 ();
 FILLCELL_X2 FILLER_0_12_86 ();
 FILLCELL_X1 FILLER_0_12_88 ();
 FILLCELL_X1 FILLER_0_12_111 ();
 FILLCELL_X4 FILLER_0_12_129 ();
 FILLCELL_X1 FILLER_0_12_133 ();
 FILLCELL_X2 FILLER_0_12_163 ();
 FILLCELL_X4 FILLER_0_12_174 ();
 FILLCELL_X1 FILLER_0_12_178 ();
 FILLCELL_X2 FILLER_0_12_186 ();
 FILLCELL_X8 FILLER_0_12_198 ();
 FILLCELL_X2 FILLER_0_12_206 ();
 FILLCELL_X1 FILLER_0_12_208 ();
 FILLCELL_X4 FILLER_0_12_225 ();
 FILLCELL_X2 FILLER_0_12_229 ();
 FILLCELL_X2 FILLER_0_12_249 ();
 FILLCELL_X1 FILLER_0_12_256 ();
 FILLCELL_X2 FILLER_0_12_261 ();
 FILLCELL_X1 FILLER_0_12_278 ();
 FILLCELL_X1 FILLER_0_12_296 ();
 FILLCELL_X2 FILLER_0_12_310 ();
 FILLCELL_X2 FILLER_0_12_316 ();
 FILLCELL_X1 FILLER_0_12_318 ();
 FILLCELL_X2 FILLER_0_12_328 ();
 FILLCELL_X1 FILLER_0_12_330 ();
 FILLCELL_X2 FILLER_0_12_334 ();
 FILLCELL_X1 FILLER_0_12_336 ();
 FILLCELL_X1 FILLER_0_12_350 ();
 FILLCELL_X1 FILLER_0_12_358 ();
 FILLCELL_X1 FILLER_0_12_365 ();
 FILLCELL_X2 FILLER_0_12_386 ();
 FILLCELL_X4 FILLER_0_13_1 ();
 FILLCELL_X2 FILLER_0_13_5 ();
 FILLCELL_X1 FILLER_0_13_7 ();
 FILLCELL_X4 FILLER_0_13_25 ();
 FILLCELL_X1 FILLER_0_13_35 ();
 FILLCELL_X1 FILLER_0_13_42 ();
 FILLCELL_X1 FILLER_0_13_53 ();
 FILLCELL_X4 FILLER_0_13_63 ();
 FILLCELL_X2 FILLER_0_13_70 ();
 FILLCELL_X1 FILLER_0_13_72 ();
 FILLCELL_X2 FILLER_0_13_89 ();
 FILLCELL_X1 FILLER_0_13_95 ();
 FILLCELL_X1 FILLER_0_13_100 ();
 FILLCELL_X1 FILLER_0_13_104 ();
 FILLCELL_X2 FILLER_0_13_115 ();
 FILLCELL_X2 FILLER_0_13_146 ();
 FILLCELL_X4 FILLER_0_13_154 ();
 FILLCELL_X1 FILLER_0_13_158 ();
 FILLCELL_X4 FILLER_0_13_171 ();
 FILLCELL_X1 FILLER_0_13_185 ();
 FILLCELL_X2 FILLER_0_13_190 ();
 FILLCELL_X2 FILLER_0_13_198 ();
 FILLCELL_X2 FILLER_0_13_206 ();
 FILLCELL_X1 FILLER_0_13_208 ();
 FILLCELL_X2 FILLER_0_13_261 ();
 FILLCELL_X2 FILLER_0_13_285 ();
 FILLCELL_X1 FILLER_0_13_296 ();
 FILLCELL_X1 FILLER_0_13_300 ();
 FILLCELL_X1 FILLER_0_13_307 ();
 FILLCELL_X1 FILLER_0_13_321 ();
 FILLCELL_X4 FILLER_0_13_326 ();
 FILLCELL_X2 FILLER_0_13_349 ();
 FILLCELL_X2 FILLER_0_13_354 ();
 FILLCELL_X2 FILLER_0_13_374 ();
 FILLCELL_X2 FILLER_0_13_379 ();
 FILLCELL_X8 FILLER_0_14_1 ();
 FILLCELL_X1 FILLER_0_14_22 ();
 FILLCELL_X1 FILLER_0_14_35 ();
 FILLCELL_X1 FILLER_0_14_46 ();
 FILLCELL_X4 FILLER_0_14_57 ();
 FILLCELL_X2 FILLER_0_14_61 ();
 FILLCELL_X8 FILLER_0_14_69 ();
 FILLCELL_X2 FILLER_0_14_77 ();
 FILLCELL_X1 FILLER_0_14_79 ();
 FILLCELL_X2 FILLER_0_14_90 ();
 FILLCELL_X1 FILLER_0_14_97 ();
 FILLCELL_X2 FILLER_0_14_114 ();
 FILLCELL_X1 FILLER_0_14_119 ();
 FILLCELL_X1 FILLER_0_14_126 ();
 FILLCELL_X1 FILLER_0_14_136 ();
 FILLCELL_X2 FILLER_0_14_169 ();
 FILLCELL_X1 FILLER_0_14_188 ();
 FILLCELL_X2 FILLER_0_14_198 ();
 FILLCELL_X1 FILLER_0_14_200 ();
 FILLCELL_X1 FILLER_0_14_228 ();
 FILLCELL_X2 FILLER_0_14_232 ();
 FILLCELL_X2 FILLER_0_14_240 ();
 FILLCELL_X2 FILLER_0_14_248 ();
 FILLCELL_X4 FILLER_0_14_263 ();
 FILLCELL_X2 FILLER_0_14_271 ();
 FILLCELL_X8 FILLER_0_14_297 ();
 FILLCELL_X4 FILLER_0_14_305 ();
 FILLCELL_X2 FILLER_0_14_309 ();
 FILLCELL_X1 FILLER_0_14_333 ();
 FILLCELL_X2 FILLER_0_14_354 ();
 FILLCELL_X1 FILLER_0_14_356 ();
 FILLCELL_X1 FILLER_0_14_377 ();
 FILLCELL_X4 FILLER_0_15_1 ();
 FILLCELL_X2 FILLER_0_15_5 ();
 FILLCELL_X1 FILLER_0_15_7 ();
 FILLCELL_X16 FILLER_0_15_15 ();
 FILLCELL_X4 FILLER_0_15_31 ();
 FILLCELL_X1 FILLER_0_15_35 ();
 FILLCELL_X2 FILLER_0_15_47 ();
 FILLCELL_X2 FILLER_0_15_55 ();
 FILLCELL_X1 FILLER_0_15_57 ();
 FILLCELL_X1 FILLER_0_15_80 ();
 FILLCELL_X8 FILLER_0_15_91 ();
 FILLCELL_X8 FILLER_0_15_105 ();
 FILLCELL_X4 FILLER_0_15_113 ();
 FILLCELL_X1 FILLER_0_15_136 ();
 FILLCELL_X1 FILLER_0_15_141 ();
 FILLCELL_X4 FILLER_0_15_146 ();
 FILLCELL_X2 FILLER_0_15_152 ();
 FILLCELL_X2 FILLER_0_15_160 ();
 FILLCELL_X2 FILLER_0_15_165 ();
 FILLCELL_X1 FILLER_0_15_177 ();
 FILLCELL_X1 FILLER_0_15_188 ();
 FILLCELL_X2 FILLER_0_15_199 ();
 FILLCELL_X2 FILLER_0_15_207 ();
 FILLCELL_X1 FILLER_0_15_209 ();
 FILLCELL_X2 FILLER_0_15_219 ();
 FILLCELL_X4 FILLER_0_15_224 ();
 FILLCELL_X1 FILLER_0_15_228 ();
 FILLCELL_X2 FILLER_0_15_239 ();
 FILLCELL_X1 FILLER_0_15_241 ();
 FILLCELL_X4 FILLER_0_15_251 ();
 FILLCELL_X1 FILLER_0_15_255 ();
 FILLCELL_X8 FILLER_0_15_269 ();
 FILLCELL_X1 FILLER_0_15_277 ();
 FILLCELL_X1 FILLER_0_15_284 ();
 FILLCELL_X4 FILLER_0_15_302 ();
 FILLCELL_X1 FILLER_0_15_306 ();
 FILLCELL_X1 FILLER_0_15_326 ();
 FILLCELL_X2 FILLER_0_15_333 ();
 FILLCELL_X1 FILLER_0_15_335 ();
 FILLCELL_X2 FILLER_0_15_342 ();
 FILLCELL_X1 FILLER_0_15_344 ();
 FILLCELL_X1 FILLER_0_15_355 ();
 FILLCELL_X16 FILLER_0_15_372 ();
 FILLCELL_X4 FILLER_0_16_1 ();
 FILLCELL_X2 FILLER_0_16_5 ();
 FILLCELL_X8 FILLER_0_16_24 ();
 FILLCELL_X8 FILLER_0_16_38 ();
 FILLCELL_X1 FILLER_0_16_46 ();
 FILLCELL_X1 FILLER_0_16_64 ();
 FILLCELL_X2 FILLER_0_16_71 ();
 FILLCELL_X1 FILLER_0_16_77 ();
 FILLCELL_X2 FILLER_0_16_84 ();
 FILLCELL_X2 FILLER_0_16_90 ();
 FILLCELL_X1 FILLER_0_16_92 ();
 FILLCELL_X4 FILLER_0_16_100 ();
 FILLCELL_X4 FILLER_0_16_107 ();
 FILLCELL_X2 FILLER_0_16_111 ();
 FILLCELL_X1 FILLER_0_16_119 ();
 FILLCELL_X1 FILLER_0_16_137 ();
 FILLCELL_X8 FILLER_0_16_148 ();
 FILLCELL_X2 FILLER_0_16_156 ();
 FILLCELL_X1 FILLER_0_16_158 ();
 FILLCELL_X1 FILLER_0_16_171 ();
 FILLCELL_X4 FILLER_0_16_175 ();
 FILLCELL_X2 FILLER_0_16_179 ();
 FILLCELL_X1 FILLER_0_16_187 ();
 FILLCELL_X1 FILLER_0_16_192 ();
 FILLCELL_X4 FILLER_0_16_197 ();
 FILLCELL_X4 FILLER_0_16_218 ();
 FILLCELL_X1 FILLER_0_16_245 ();
 FILLCELL_X2 FILLER_0_16_254 ();
 FILLCELL_X2 FILLER_0_16_262 ();
 FILLCELL_X2 FILLER_0_16_289 ();
 FILLCELL_X1 FILLER_0_16_291 ();
 FILLCELL_X1 FILLER_0_16_309 ();
 FILLCELL_X1 FILLER_0_16_314 ();
 FILLCELL_X1 FILLER_0_16_317 ();
 FILLCELL_X1 FILLER_0_16_336 ();
 FILLCELL_X1 FILLER_0_16_340 ();
 FILLCELL_X1 FILLER_0_16_347 ();
 FILLCELL_X1 FILLER_0_16_351 ();
 FILLCELL_X2 FILLER_0_16_358 ();
 FILLCELL_X8 FILLER_0_16_380 ();
 FILLCELL_X16 FILLER_0_17_1 ();
 FILLCELL_X4 FILLER_0_17_17 ();
 FILLCELL_X2 FILLER_0_17_21 ();
 FILLCELL_X4 FILLER_0_17_40 ();
 FILLCELL_X1 FILLER_0_17_44 ();
 FILLCELL_X2 FILLER_0_17_51 ();
 FILLCELL_X1 FILLER_0_17_53 ();
 FILLCELL_X4 FILLER_0_17_60 ();
 FILLCELL_X1 FILLER_0_17_64 ();
 FILLCELL_X1 FILLER_0_17_71 ();
 FILLCELL_X1 FILLER_0_17_78 ();
 FILLCELL_X2 FILLER_0_17_83 ();
 FILLCELL_X4 FILLER_0_17_101 ();
 FILLCELL_X2 FILLER_0_17_105 ();
 FILLCELL_X1 FILLER_0_17_107 ();
 FILLCELL_X2 FILLER_0_17_131 ();
 FILLCELL_X1 FILLER_0_17_137 ();
 FILLCELL_X4 FILLER_0_17_158 ();
 FILLCELL_X1 FILLER_0_17_177 ();
 FILLCELL_X2 FILLER_0_17_196 ();
 FILLCELL_X1 FILLER_0_17_204 ();
 FILLCELL_X4 FILLER_0_17_208 ();
 FILLCELL_X2 FILLER_0_17_212 ();
 FILLCELL_X1 FILLER_0_17_214 ();
 FILLCELL_X16 FILLER_0_17_218 ();
 FILLCELL_X1 FILLER_0_17_234 ();
 FILLCELL_X1 FILLER_0_17_246 ();
 FILLCELL_X4 FILLER_0_17_251 ();
 FILLCELL_X1 FILLER_0_17_255 ();
 FILLCELL_X1 FILLER_0_17_269 ();
 FILLCELL_X1 FILLER_0_17_276 ();
 FILLCELL_X1 FILLER_0_17_280 ();
 FILLCELL_X8 FILLER_0_17_294 ();
 FILLCELL_X1 FILLER_0_17_326 ();
 FILLCELL_X2 FILLER_0_17_331 ();
 FILLCELL_X2 FILLER_0_17_344 ();
 FILLCELL_X2 FILLER_0_17_357 ();
 FILLCELL_X2 FILLER_0_17_386 ();
 FILLCELL_X16 FILLER_0_18_1 ();
 FILLCELL_X2 FILLER_0_18_17 ();
 FILLCELL_X1 FILLER_0_18_19 ();
 FILLCELL_X1 FILLER_0_18_26 ();
 FILLCELL_X2 FILLER_0_18_44 ();
 FILLCELL_X1 FILLER_0_18_70 ();
 FILLCELL_X8 FILLER_0_18_80 ();
 FILLCELL_X1 FILLER_0_18_88 ();
 FILLCELL_X4 FILLER_0_18_90 ();
 FILLCELL_X2 FILLER_0_18_94 ();
 FILLCELL_X1 FILLER_0_18_117 ();
 FILLCELL_X2 FILLER_0_18_156 ();
 FILLCELL_X4 FILLER_0_18_167 ();
 FILLCELL_X1 FILLER_0_18_171 ();
 FILLCELL_X4 FILLER_0_18_188 ();
 FILLCELL_X4 FILLER_0_18_201 ();
 FILLCELL_X2 FILLER_0_18_254 ();
 FILLCELL_X1 FILLER_0_18_260 ();
 FILLCELL_X1 FILLER_0_18_268 ();
 FILLCELL_X1 FILLER_0_18_273 ();
 FILLCELL_X1 FILLER_0_18_278 ();
 FILLCELL_X1 FILLER_0_18_285 ();
 FILLCELL_X2 FILLER_0_18_293 ();
 FILLCELL_X1 FILLER_0_18_295 ();
 FILLCELL_X1 FILLER_0_18_307 ();
 FILLCELL_X2 FILLER_0_18_316 ();
 FILLCELL_X1 FILLER_0_18_318 ();
 FILLCELL_X4 FILLER_0_18_336 ();
 FILLCELL_X1 FILLER_0_18_340 ();
 FILLCELL_X1 FILLER_0_18_347 ();
 FILLCELL_X2 FILLER_0_18_350 ();
 FILLCELL_X2 FILLER_0_18_356 ();
 FILLCELL_X1 FILLER_0_18_358 ();
 FILLCELL_X2 FILLER_0_18_365 ();
 FILLCELL_X1 FILLER_0_18_367 ();
 FILLCELL_X2 FILLER_0_18_372 ();
 FILLCELL_X2 FILLER_0_18_382 ();
 FILLCELL_X1 FILLER_0_18_387 ();
 FILLCELL_X16 FILLER_0_19_1 ();
 FILLCELL_X1 FILLER_0_19_17 ();
 FILLCELL_X1 FILLER_0_19_22 ();
 FILLCELL_X4 FILLER_0_19_27 ();
 FILLCELL_X2 FILLER_0_19_31 ();
 FILLCELL_X1 FILLER_0_19_33 ();
 FILLCELL_X1 FILLER_0_19_55 ();
 FILLCELL_X1 FILLER_0_19_59 ();
 FILLCELL_X1 FILLER_0_19_69 ();
 FILLCELL_X2 FILLER_0_19_80 ();
 FILLCELL_X1 FILLER_0_19_82 ();
 FILLCELL_X1 FILLER_0_19_96 ();
 FILLCELL_X1 FILLER_0_19_101 ();
 FILLCELL_X1 FILLER_0_19_105 ();
 FILLCELL_X1 FILLER_0_19_111 ();
 FILLCELL_X2 FILLER_0_19_115 ();
 FILLCELL_X1 FILLER_0_19_121 ();
 FILLCELL_X2 FILLER_0_19_128 ();
 FILLCELL_X1 FILLER_0_19_130 ();
 FILLCELL_X4 FILLER_0_19_135 ();
 FILLCELL_X4 FILLER_0_19_142 ();
 FILLCELL_X2 FILLER_0_19_146 ();
 FILLCELL_X1 FILLER_0_19_148 ();
 FILLCELL_X4 FILLER_0_19_155 ();
 FILLCELL_X2 FILLER_0_19_159 ();
 FILLCELL_X1 FILLER_0_19_161 ();
 FILLCELL_X4 FILLER_0_19_167 ();
 FILLCELL_X1 FILLER_0_19_171 ();
 FILLCELL_X8 FILLER_0_19_179 ();
 FILLCELL_X2 FILLER_0_19_187 ();
 FILLCELL_X1 FILLER_0_19_195 ();
 FILLCELL_X2 FILLER_0_19_200 ();
 FILLCELL_X4 FILLER_0_19_208 ();
 FILLCELL_X2 FILLER_0_19_212 ();
 FILLCELL_X2 FILLER_0_19_224 ();
 FILLCELL_X2 FILLER_0_19_229 ();
 FILLCELL_X4 FILLER_0_19_281 ();
 FILLCELL_X2 FILLER_0_19_285 ();
 FILLCELL_X4 FILLER_0_19_305 ();
 FILLCELL_X2 FILLER_0_19_309 ();
 FILLCELL_X4 FILLER_0_19_317 ();
 FILLCELL_X2 FILLER_0_19_333 ();
 FILLCELL_X2 FILLER_0_19_357 ();
 FILLCELL_X1 FILLER_0_19_359 ();
 FILLCELL_X8 FILLER_0_19_362 ();
 FILLCELL_X4 FILLER_0_19_373 ();
 FILLCELL_X4 FILLER_0_19_384 ();
 FILLCELL_X32 FILLER_0_20_1 ();
 FILLCELL_X2 FILLER_0_20_33 ();
 FILLCELL_X1 FILLER_0_20_35 ();
 FILLCELL_X4 FILLER_0_20_39 ();
 FILLCELL_X2 FILLER_0_20_43 ();
 FILLCELL_X1 FILLER_0_20_54 ();
 FILLCELL_X1 FILLER_0_20_65 ();
 FILLCELL_X2 FILLER_0_20_83 ();
 FILLCELL_X1 FILLER_0_20_88 ();
 FILLCELL_X1 FILLER_0_20_126 ();
 FILLCELL_X1 FILLER_0_20_133 ();
 FILLCELL_X1 FILLER_0_20_144 ();
 FILLCELL_X2 FILLER_0_20_158 ();
 FILLCELL_X1 FILLER_0_20_166 ();
 FILLCELL_X1 FILLER_0_20_169 ();
 FILLCELL_X1 FILLER_0_20_175 ();
 FILLCELL_X2 FILLER_0_20_186 ();
 FILLCELL_X1 FILLER_0_20_188 ();
 FILLCELL_X2 FILLER_0_20_229 ();
 FILLCELL_X8 FILLER_0_20_237 ();
 FILLCELL_X2 FILLER_0_20_245 ();
 FILLCELL_X1 FILLER_0_20_260 ();
 FILLCELL_X1 FILLER_0_20_266 ();
 FILLCELL_X1 FILLER_0_20_268 ();
 FILLCELL_X1 FILLER_0_20_275 ();
 FILLCELL_X1 FILLER_0_20_282 ();
 FILLCELL_X2 FILLER_0_20_302 ();
 FILLCELL_X8 FILLER_0_20_313 ();
 FILLCELL_X4 FILLER_0_20_321 ();
 FILLCELL_X1 FILLER_0_20_325 ();
 FILLCELL_X4 FILLER_0_20_358 ();
 FILLCELL_X1 FILLER_0_20_362 ();
 FILLCELL_X1 FILLER_0_20_367 ();
 FILLCELL_X1 FILLER_0_20_381 ();
 FILLCELL_X2 FILLER_0_20_385 ();
 FILLCELL_X1 FILLER_0_20_387 ();
 FILLCELL_X4 FILLER_0_21_1 ();
 FILLCELL_X4 FILLER_0_21_22 ();
 FILLCELL_X2 FILLER_0_21_54 ();
 FILLCELL_X2 FILLER_0_21_62 ();
 FILLCELL_X1 FILLER_0_21_64 ();
 FILLCELL_X2 FILLER_0_21_71 ();
 FILLCELL_X1 FILLER_0_21_73 ();
 FILLCELL_X2 FILLER_0_21_80 ();
 FILLCELL_X2 FILLER_0_21_86 ();
 FILLCELL_X1 FILLER_0_21_88 ();
 FILLCELL_X1 FILLER_0_21_108 ();
 FILLCELL_X1 FILLER_0_21_115 ();
 FILLCELL_X1 FILLER_0_21_126 ();
 FILLCELL_X4 FILLER_0_21_152 ();
 FILLCELL_X4 FILLER_0_21_162 ();
 FILLCELL_X2 FILLER_0_21_166 ();
 FILLCELL_X1 FILLER_0_21_168 ();
 FILLCELL_X2 FILLER_0_21_176 ();
 FILLCELL_X2 FILLER_0_21_185 ();
 FILLCELL_X1 FILLER_0_21_197 ();
 FILLCELL_X4 FILLER_0_21_208 ();
 FILLCELL_X2 FILLER_0_21_234 ();
 FILLCELL_X1 FILLER_0_21_236 ();
 FILLCELL_X4 FILLER_0_21_243 ();
 FILLCELL_X2 FILLER_0_21_247 ();
 FILLCELL_X1 FILLER_0_21_249 ();
 FILLCELL_X1 FILLER_0_21_268 ();
 FILLCELL_X4 FILLER_0_21_291 ();
 FILLCELL_X2 FILLER_0_21_295 ();
 FILLCELL_X4 FILLER_0_21_312 ();
 FILLCELL_X2 FILLER_0_21_316 ();
 FILLCELL_X2 FILLER_0_21_337 ();
 FILLCELL_X1 FILLER_0_21_355 ();
 FILLCELL_X2 FILLER_0_21_386 ();
 FILLCELL_X8 FILLER_0_22_1 ();
 FILLCELL_X2 FILLER_0_22_9 ();
 FILLCELL_X1 FILLER_0_22_11 ();
 FILLCELL_X2 FILLER_0_22_23 ();
 FILLCELL_X2 FILLER_0_22_27 ();
 FILLCELL_X1 FILLER_0_22_29 ();
 FILLCELL_X1 FILLER_0_22_37 ();
 FILLCELL_X4 FILLER_0_22_47 ();
 FILLCELL_X1 FILLER_0_22_51 ();
 FILLCELL_X8 FILLER_0_22_62 ();
 FILLCELL_X1 FILLER_0_22_70 ();
 FILLCELL_X2 FILLER_0_22_86 ();
 FILLCELL_X1 FILLER_0_22_88 ();
 FILLCELL_X4 FILLER_0_22_103 ();
 FILLCELL_X1 FILLER_0_22_130 ();
 FILLCELL_X1 FILLER_0_22_144 ();
 FILLCELL_X2 FILLER_0_22_148 ();
 FILLCELL_X2 FILLER_0_22_172 ();
 FILLCELL_X2 FILLER_0_22_180 ();
 FILLCELL_X1 FILLER_0_22_182 ();
 FILLCELL_X2 FILLER_0_22_195 ();
 FILLCELL_X1 FILLER_0_22_201 ();
 FILLCELL_X2 FILLER_0_22_249 ();
 FILLCELL_X2 FILLER_0_22_265 ();
 FILLCELL_X1 FILLER_0_22_268 ();
 FILLCELL_X2 FILLER_0_22_273 ();
 FILLCELL_X2 FILLER_0_22_277 ();
 FILLCELL_X2 FILLER_0_22_282 ();
 FILLCELL_X4 FILLER_0_22_302 ();
 FILLCELL_X1 FILLER_0_22_310 ();
 FILLCELL_X1 FILLER_0_22_317 ();
 FILLCELL_X1 FILLER_0_22_322 ();
 FILLCELL_X1 FILLER_0_22_329 ();
 FILLCELL_X1 FILLER_0_22_337 ();
 FILLCELL_X1 FILLER_0_22_346 ();
 FILLCELL_X8 FILLER_0_22_350 ();
 FILLCELL_X2 FILLER_0_22_358 ();
 FILLCELL_X1 FILLER_0_22_383 ();
 FILLCELL_X2 FILLER_0_23_1 ();
 FILLCELL_X1 FILLER_0_23_3 ();
 FILLCELL_X2 FILLER_0_23_27 ();
 FILLCELL_X1 FILLER_0_23_39 ();
 FILLCELL_X1 FILLER_0_23_46 ();
 FILLCELL_X1 FILLER_0_23_53 ();
 FILLCELL_X1 FILLER_0_23_63 ();
 FILLCELL_X2 FILLER_0_23_70 ();
 FILLCELL_X1 FILLER_0_23_78 ();
 FILLCELL_X1 FILLER_0_23_86 ();
 FILLCELL_X1 FILLER_0_23_93 ();
 FILLCELL_X1 FILLER_0_23_131 ();
 FILLCELL_X1 FILLER_0_23_138 ();
 FILLCELL_X1 FILLER_0_23_142 ();
 FILLCELL_X1 FILLER_0_23_149 ();
 FILLCELL_X2 FILLER_0_23_170 ();
 FILLCELL_X2 FILLER_0_23_185 ();
 FILLCELL_X2 FILLER_0_23_210 ();
 FILLCELL_X1 FILLER_0_23_212 ();
 FILLCELL_X2 FILLER_0_23_239 ();
 FILLCELL_X2 FILLER_0_23_244 ();
 FILLCELL_X2 FILLER_0_23_255 ();
 FILLCELL_X1 FILLER_0_23_257 ();
 FILLCELL_X1 FILLER_0_23_262 ();
 FILLCELL_X2 FILLER_0_23_269 ();
 FILLCELL_X2 FILLER_0_23_298 ();
 FILLCELL_X1 FILLER_0_23_300 ();
 FILLCELL_X1 FILLER_0_23_307 ();
 FILLCELL_X1 FILLER_0_23_314 ();
 FILLCELL_X4 FILLER_0_23_328 ();
 FILLCELL_X1 FILLER_0_23_332 ();
 FILLCELL_X4 FILLER_0_23_339 ();
 FILLCELL_X4 FILLER_0_23_352 ();
 FILLCELL_X1 FILLER_0_23_363 ();
 FILLCELL_X1 FILLER_0_23_383 ();
 FILLCELL_X2 FILLER_0_23_386 ();
 FILLCELL_X4 FILLER_0_24_1 ();
 FILLCELL_X1 FILLER_0_24_5 ();
 FILLCELL_X8 FILLER_0_24_17 ();
 FILLCELL_X2 FILLER_0_24_25 ();
 FILLCELL_X1 FILLER_0_24_27 ();
 FILLCELL_X2 FILLER_0_24_37 ();
 FILLCELL_X1 FILLER_0_24_54 ();
 FILLCELL_X8 FILLER_0_24_66 ();
 FILLCELL_X2 FILLER_0_24_74 ();
 FILLCELL_X1 FILLER_0_24_76 ();
 FILLCELL_X1 FILLER_0_24_88 ();
 FILLCELL_X4 FILLER_0_24_96 ();
 FILLCELL_X2 FILLER_0_24_100 ();
 FILLCELL_X1 FILLER_0_24_102 ();
 FILLCELL_X1 FILLER_0_24_118 ();
 FILLCELL_X2 FILLER_0_24_143 ();
 FILLCELL_X1 FILLER_0_24_151 ();
 FILLCELL_X1 FILLER_0_24_158 ();
 FILLCELL_X1 FILLER_0_24_163 ();
 FILLCELL_X2 FILLER_0_24_168 ();
 FILLCELL_X2 FILLER_0_24_173 ();
 FILLCELL_X1 FILLER_0_24_175 ();
 FILLCELL_X2 FILLER_0_24_197 ();
 FILLCELL_X2 FILLER_0_24_249 ();
 FILLCELL_X1 FILLER_0_24_257 ();
 FILLCELL_X2 FILLER_0_24_264 ();
 FILLCELL_X1 FILLER_0_24_266 ();
 FILLCELL_X1 FILLER_0_24_268 ();
 FILLCELL_X1 FILLER_0_24_286 ();
 FILLCELL_X1 FILLER_0_24_290 ();
 FILLCELL_X1 FILLER_0_24_300 ();
 FILLCELL_X4 FILLER_0_24_314 ();
 FILLCELL_X2 FILLER_0_24_328 ();
 FILLCELL_X1 FILLER_0_24_330 ();
 FILLCELL_X4 FILLER_0_24_340 ();
 FILLCELL_X1 FILLER_0_24_362 ();
 FILLCELL_X1 FILLER_0_24_367 ();
 FILLCELL_X1 FILLER_0_24_370 ();
 FILLCELL_X1 FILLER_0_24_380 ();
 FILLCELL_X1 FILLER_0_24_387 ();
 FILLCELL_X4 FILLER_0_25_25 ();
 FILLCELL_X2 FILLER_0_25_29 ();
 FILLCELL_X1 FILLER_0_25_31 ();
 FILLCELL_X4 FILLER_0_25_36 ();
 FILLCELL_X1 FILLER_0_25_46 ();
 FILLCELL_X2 FILLER_0_25_70 ();
 FILLCELL_X4 FILLER_0_25_88 ();
 FILLCELL_X4 FILLER_0_25_106 ();
 FILLCELL_X2 FILLER_0_25_110 ();
 FILLCELL_X1 FILLER_0_25_112 ();
 FILLCELL_X2 FILLER_0_25_116 ();
 FILLCELL_X1 FILLER_0_25_124 ();
 FILLCELL_X2 FILLER_0_25_135 ();
 FILLCELL_X1 FILLER_0_25_137 ();
 FILLCELL_X1 FILLER_0_25_144 ();
 FILLCELL_X1 FILLER_0_25_159 ();
 FILLCELL_X1 FILLER_0_25_163 ();
 FILLCELL_X1 FILLER_0_25_170 ();
 FILLCELL_X1 FILLER_0_25_174 ();
 FILLCELL_X4 FILLER_0_25_197 ();
 FILLCELL_X2 FILLER_0_25_201 ();
 FILLCELL_X1 FILLER_0_25_203 ();
 FILLCELL_X2 FILLER_0_25_207 ();
 FILLCELL_X1 FILLER_0_25_209 ();
 FILLCELL_X1 FILLER_0_25_214 ();
 FILLCELL_X8 FILLER_0_25_260 ();
 FILLCELL_X2 FILLER_0_25_268 ();
 FILLCELL_X16 FILLER_0_25_280 ();
 FILLCELL_X8 FILLER_0_25_296 ();
 FILLCELL_X2 FILLER_0_25_304 ();
 FILLCELL_X2 FILLER_0_25_326 ();
 FILLCELL_X8 FILLER_0_25_334 ();
 FILLCELL_X2 FILLER_0_25_342 ();
 FILLCELL_X1 FILLER_0_25_344 ();
 FILLCELL_X1 FILLER_0_25_355 ();
 FILLCELL_X2 FILLER_0_25_360 ();
 FILLCELL_X1 FILLER_0_25_381 ();
 FILLCELL_X2 FILLER_0_25_385 ();
 FILLCELL_X1 FILLER_0_25_387 ();
 FILLCELL_X2 FILLER_0_26_25 ();
 FILLCELL_X1 FILLER_0_26_27 ();
 FILLCELL_X2 FILLER_0_26_37 ();
 FILLCELL_X1 FILLER_0_26_39 ();
 FILLCELL_X1 FILLER_0_26_49 ();
 FILLCELL_X4 FILLER_0_26_62 ();
 FILLCELL_X4 FILLER_0_26_69 ();
 FILLCELL_X1 FILLER_0_26_90 ();
 FILLCELL_X1 FILLER_0_26_102 ();
 FILLCELL_X1 FILLER_0_26_112 ();
 FILLCELL_X1 FILLER_0_26_116 ();
 FILLCELL_X1 FILLER_0_26_123 ();
 FILLCELL_X1 FILLER_0_26_136 ();
 FILLCELL_X1 FILLER_0_26_140 ();
 FILLCELL_X1 FILLER_0_26_143 ();
 FILLCELL_X4 FILLER_0_26_158 ();
 FILLCELL_X2 FILLER_0_26_162 ();
 FILLCELL_X4 FILLER_0_26_172 ();
 FILLCELL_X2 FILLER_0_26_193 ();
 FILLCELL_X4 FILLER_0_26_233 ();
 FILLCELL_X2 FILLER_0_26_237 ();
 FILLCELL_X1 FILLER_0_26_239 ();
 FILLCELL_X8 FILLER_0_26_244 ();
 FILLCELL_X2 FILLER_0_26_252 ();
 FILLCELL_X1 FILLER_0_26_254 ();
 FILLCELL_X2 FILLER_0_26_265 ();
 FILLCELL_X2 FILLER_0_26_268 ();
 FILLCELL_X1 FILLER_0_26_270 ();
 FILLCELL_X2 FILLER_0_26_290 ();
 FILLCELL_X1 FILLER_0_26_292 ();
 FILLCELL_X2 FILLER_0_26_305 ();
 FILLCELL_X8 FILLER_0_26_312 ();
 FILLCELL_X1 FILLER_0_26_320 ();
 FILLCELL_X2 FILLER_0_26_332 ();
 FILLCELL_X1 FILLER_0_26_334 ();
 FILLCELL_X8 FILLER_0_26_345 ();
 FILLCELL_X1 FILLER_0_26_355 ();
 FILLCELL_X1 FILLER_0_26_360 ();
 FILLCELL_X1 FILLER_0_26_367 ();
 FILLCELL_X2 FILLER_0_26_374 ();
 FILLCELL_X8 FILLER_0_26_380 ();
 FILLCELL_X1 FILLER_0_27_1 ();
 FILLCELL_X1 FILLER_0_27_6 ();
 FILLCELL_X1 FILLER_0_27_13 ();
 FILLCELL_X1 FILLER_0_27_17 ();
 FILLCELL_X1 FILLER_0_27_24 ();
 FILLCELL_X2 FILLER_0_27_34 ();
 FILLCELL_X1 FILLER_0_27_36 ();
 FILLCELL_X1 FILLER_0_27_46 ();
 FILLCELL_X2 FILLER_0_27_54 ();
 FILLCELL_X1 FILLER_0_27_65 ();
 FILLCELL_X1 FILLER_0_27_75 ();
 FILLCELL_X2 FILLER_0_27_87 ();
 FILLCELL_X4 FILLER_0_27_122 ();
 FILLCELL_X2 FILLER_0_27_126 ();
 FILLCELL_X8 FILLER_0_27_134 ();
 FILLCELL_X2 FILLER_0_27_142 ();
 FILLCELL_X1 FILLER_0_27_144 ();
 FILLCELL_X2 FILLER_0_27_151 ();
 FILLCELL_X1 FILLER_0_27_159 ();
 FILLCELL_X2 FILLER_0_27_166 ();
 FILLCELL_X1 FILLER_0_27_168 ();
 FILLCELL_X4 FILLER_0_27_182 ();
 FILLCELL_X2 FILLER_0_27_186 ();
 FILLCELL_X1 FILLER_0_27_188 ();
 FILLCELL_X2 FILLER_0_27_208 ();
 FILLCELL_X2 FILLER_0_27_213 ();
 FILLCELL_X1 FILLER_0_27_215 ();
 FILLCELL_X8 FILLER_0_27_222 ();
 FILLCELL_X1 FILLER_0_27_230 ();
 FILLCELL_X2 FILLER_0_27_253 ();
 FILLCELL_X2 FILLER_0_27_270 ();
 FILLCELL_X4 FILLER_0_27_274 ();
 FILLCELL_X8 FILLER_0_27_299 ();
 FILLCELL_X4 FILLER_0_27_307 ();
 FILLCELL_X1 FILLER_0_27_311 ();
 FILLCELL_X8 FILLER_0_27_322 ();
 FILLCELL_X2 FILLER_0_27_330 ();
 FILLCELL_X4 FILLER_0_27_342 ();
 FILLCELL_X1 FILLER_0_27_346 ();
 FILLCELL_X8 FILLER_0_27_357 ();
 FILLCELL_X4 FILLER_0_27_365 ();
 FILLCELL_X2 FILLER_0_27_369 ();
 FILLCELL_X4 FILLER_0_28_1 ();
 FILLCELL_X1 FILLER_0_28_5 ();
 FILLCELL_X1 FILLER_0_28_12 ();
 FILLCELL_X1 FILLER_0_28_17 ();
 FILLCELL_X8 FILLER_0_28_21 ();
 FILLCELL_X1 FILLER_0_28_29 ();
 FILLCELL_X4 FILLER_0_28_36 ();
 FILLCELL_X1 FILLER_0_28_99 ();
 FILLCELL_X2 FILLER_0_28_106 ();
 FILLCELL_X1 FILLER_0_28_108 ();
 FILLCELL_X1 FILLER_0_28_131 ();
 FILLCELL_X2 FILLER_0_28_136 ();
 FILLCELL_X1 FILLER_0_28_142 ();
 FILLCELL_X2 FILLER_0_28_149 ();
 FILLCELL_X2 FILLER_0_28_154 ();
 FILLCELL_X2 FILLER_0_28_162 ();
 FILLCELL_X1 FILLER_0_28_193 ();
 FILLCELL_X2 FILLER_0_28_196 ();
 FILLCELL_X2 FILLER_0_28_201 ();
 FILLCELL_X4 FILLER_0_28_209 ();
 FILLCELL_X2 FILLER_0_28_226 ();
 FILLCELL_X4 FILLER_0_28_231 ();
 FILLCELL_X1 FILLER_0_28_250 ();
 FILLCELL_X1 FILLER_0_28_255 ();
 FILLCELL_X1 FILLER_0_28_262 ();
 FILLCELL_X8 FILLER_0_28_303 ();
 FILLCELL_X2 FILLER_0_28_311 ();
 FILLCELL_X1 FILLER_0_28_343 ();
 FILLCELL_X2 FILLER_0_28_361 ();
 FILLCELL_X8 FILLER_0_29_1 ();
 FILLCELL_X1 FILLER_0_29_13 ();
 FILLCELL_X1 FILLER_0_29_18 ();
 FILLCELL_X2 FILLER_0_29_25 ();
 FILLCELL_X1 FILLER_0_29_27 ();
 FILLCELL_X2 FILLER_0_29_38 ();
 FILLCELL_X2 FILLER_0_29_44 ();
 FILLCELL_X2 FILLER_0_29_56 ();
 FILLCELL_X1 FILLER_0_29_87 ();
 FILLCELL_X1 FILLER_0_29_93 ();
 FILLCELL_X2 FILLER_0_29_106 ();
 FILLCELL_X1 FILLER_0_29_108 ();
 FILLCELL_X8 FILLER_0_29_113 ();
 FILLCELL_X2 FILLER_0_29_127 ();
 FILLCELL_X1 FILLER_0_29_129 ();
 FILLCELL_X4 FILLER_0_29_163 ();
 FILLCELL_X1 FILLER_0_29_167 ();
 FILLCELL_X2 FILLER_0_29_174 ();
 FILLCELL_X8 FILLER_0_29_182 ();
 FILLCELL_X1 FILLER_0_29_203 ();
 FILLCELL_X1 FILLER_0_29_224 ();
 FILLCELL_X2 FILLER_0_29_242 ();
 FILLCELL_X1 FILLER_0_29_247 ();
 FILLCELL_X2 FILLER_0_29_254 ();
 FILLCELL_X2 FILLER_0_29_260 ();
 FILLCELL_X2 FILLER_0_29_287 ();
 FILLCELL_X2 FILLER_0_29_291 ();
 FILLCELL_X1 FILLER_0_29_293 ();
 FILLCELL_X4 FILLER_0_29_306 ();
 FILLCELL_X1 FILLER_0_29_310 ();
 FILLCELL_X2 FILLER_0_29_317 ();
 FILLCELL_X2 FILLER_0_29_325 ();
 FILLCELL_X1 FILLER_0_29_357 ();
 FILLCELL_X1 FILLER_0_29_361 ();
 FILLCELL_X1 FILLER_0_29_365 ();
 FILLCELL_X1 FILLER_0_29_372 ();
 FILLCELL_X1 FILLER_0_29_384 ();
 FILLCELL_X4 FILLER_0_30_1 ();
 FILLCELL_X2 FILLER_0_30_5 ();
 FILLCELL_X1 FILLER_0_30_32 ();
 FILLCELL_X1 FILLER_0_30_36 ();
 FILLCELL_X1 FILLER_0_30_43 ();
 FILLCELL_X1 FILLER_0_30_50 ();
 FILLCELL_X1 FILLER_0_30_65 ();
 FILLCELL_X8 FILLER_0_30_72 ();
 FILLCELL_X2 FILLER_0_30_83 ();
 FILLCELL_X1 FILLER_0_30_85 ();
 FILLCELL_X1 FILLER_0_30_90 ();
 FILLCELL_X4 FILLER_0_30_101 ();
 FILLCELL_X4 FILLER_0_30_108 ();
 FILLCELL_X4 FILLER_0_30_122 ();
 FILLCELL_X2 FILLER_0_30_126 ();
 FILLCELL_X1 FILLER_0_30_128 ();
 FILLCELL_X2 FILLER_0_30_135 ();
 FILLCELL_X4 FILLER_0_30_149 ();
 FILLCELL_X1 FILLER_0_30_173 ();
 FILLCELL_X4 FILLER_0_30_178 ();
 FILLCELL_X4 FILLER_0_30_199 ();
 FILLCELL_X1 FILLER_0_30_203 ();
 FILLCELL_X2 FILLER_0_30_214 ();
 FILLCELL_X1 FILLER_0_30_216 ();
 FILLCELL_X2 FILLER_0_30_249 ();
 FILLCELL_X4 FILLER_0_30_261 ();
 FILLCELL_X2 FILLER_0_30_265 ();
 FILLCELL_X1 FILLER_0_30_268 ();
 FILLCELL_X1 FILLER_0_30_281 ();
 FILLCELL_X2 FILLER_0_30_286 ();
 FILLCELL_X2 FILLER_0_30_294 ();
 FILLCELL_X2 FILLER_0_30_300 ();
 FILLCELL_X1 FILLER_0_30_302 ();
 FILLCELL_X2 FILLER_0_30_324 ();
 FILLCELL_X1 FILLER_0_30_339 ();
 FILLCELL_X1 FILLER_0_30_346 ();
 FILLCELL_X2 FILLER_0_30_350 ();
 FILLCELL_X1 FILLER_0_30_358 ();
 FILLCELL_X2 FILLER_0_30_362 ();
 FILLCELL_X1 FILLER_0_30_370 ();
 FILLCELL_X4 FILLER_0_30_384 ();
 FILLCELL_X4 FILLER_0_31_1 ();
 FILLCELL_X2 FILLER_0_31_5 ();
 FILLCELL_X1 FILLER_0_31_24 ();
 FILLCELL_X2 FILLER_0_31_43 ();
 FILLCELL_X2 FILLER_0_31_48 ();
 FILLCELL_X2 FILLER_0_31_53 ();
 FILLCELL_X1 FILLER_0_31_55 ();
 FILLCELL_X4 FILLER_0_31_62 ();
 FILLCELL_X2 FILLER_0_31_66 ();
 FILLCELL_X1 FILLER_0_31_68 ();
 FILLCELL_X4 FILLER_0_31_77 ();
 FILLCELL_X1 FILLER_0_31_81 ();
 FILLCELL_X4 FILLER_0_31_85 ();
 FILLCELL_X2 FILLER_0_31_89 ();
 FILLCELL_X1 FILLER_0_31_91 ();
 FILLCELL_X2 FILLER_0_31_119 ();
 FILLCELL_X8 FILLER_0_31_141 ();
 FILLCELL_X4 FILLER_0_31_149 ();
 FILLCELL_X2 FILLER_0_31_153 ();
 FILLCELL_X1 FILLER_0_31_155 ();
 FILLCELL_X4 FILLER_0_31_165 ();
 FILLCELL_X2 FILLER_0_31_169 ();
 FILLCELL_X1 FILLER_0_31_171 ();
 FILLCELL_X4 FILLER_0_31_179 ();
 FILLCELL_X2 FILLER_0_31_183 ();
 FILLCELL_X1 FILLER_0_31_185 ();
 FILLCELL_X2 FILLER_0_31_192 ();
 FILLCELL_X4 FILLER_0_31_200 ();
 FILLCELL_X2 FILLER_0_31_204 ();
 FILLCELL_X4 FILLER_0_31_227 ();
 FILLCELL_X1 FILLER_0_31_259 ();
 FILLCELL_X1 FILLER_0_31_266 ();
 FILLCELL_X1 FILLER_0_31_276 ();
 FILLCELL_X1 FILLER_0_31_281 ();
 FILLCELL_X2 FILLER_0_31_292 ();
 FILLCELL_X1 FILLER_0_31_294 ();
 FILLCELL_X2 FILLER_0_31_301 ();
 FILLCELL_X1 FILLER_0_31_303 ();
 FILLCELL_X2 FILLER_0_31_323 ();
 FILLCELL_X2 FILLER_0_31_332 ();
 FILLCELL_X2 FILLER_0_31_344 ();
 FILLCELL_X1 FILLER_0_31_355 ();
 FILLCELL_X1 FILLER_0_31_366 ();
 FILLCELL_X2 FILLER_0_31_370 ();
 FILLCELL_X4 FILLER_0_31_384 ();
 FILLCELL_X1 FILLER_0_32_33 ();
 FILLCELL_X8 FILLER_0_32_60 ();
 FILLCELL_X2 FILLER_0_32_68 ();
 FILLCELL_X1 FILLER_0_32_70 ();
 FILLCELL_X1 FILLER_0_32_82 ();
 FILLCELL_X8 FILLER_0_32_93 ();
 FILLCELL_X2 FILLER_0_32_111 ();
 FILLCELL_X1 FILLER_0_32_155 ();
 FILLCELL_X4 FILLER_0_32_170 ();
 FILLCELL_X2 FILLER_0_32_174 ();
 FILLCELL_X1 FILLER_0_32_176 ();
 FILLCELL_X2 FILLER_0_32_190 ();
 FILLCELL_X1 FILLER_0_32_192 ();
 FILLCELL_X4 FILLER_0_32_201 ();
 FILLCELL_X1 FILLER_0_32_205 ();
 FILLCELL_X1 FILLER_0_32_215 ();
 FILLCELL_X1 FILLER_0_32_260 ();
 FILLCELL_X1 FILLER_0_32_284 ();
 FILLCELL_X2 FILLER_0_32_289 ();
 FILLCELL_X1 FILLER_0_32_291 ();
 FILLCELL_X2 FILLER_0_32_302 ();
 FILLCELL_X4 FILLER_0_32_308 ();
 FILLCELL_X1 FILLER_0_32_324 ();
 FILLCELL_X8 FILLER_0_32_331 ();
 FILLCELL_X2 FILLER_0_32_339 ();
 FILLCELL_X1 FILLER_0_32_350 ();
 FILLCELL_X1 FILLER_0_32_364 ();
 FILLCELL_X1 FILLER_0_32_369 ();
 FILLCELL_X8 FILLER_0_32_380 ();
 FILLCELL_X8 FILLER_0_33_1 ();
 FILLCELL_X1 FILLER_0_33_17 ();
 FILLCELL_X1 FILLER_0_33_29 ();
 FILLCELL_X1 FILLER_0_33_36 ();
 FILLCELL_X2 FILLER_0_33_41 ();
 FILLCELL_X2 FILLER_0_33_46 ();
 FILLCELL_X2 FILLER_0_33_54 ();
 FILLCELL_X4 FILLER_0_33_59 ();
 FILLCELL_X2 FILLER_0_33_101 ();
 FILLCELL_X1 FILLER_0_33_120 ();
 FILLCELL_X1 FILLER_0_33_127 ();
 FILLCELL_X1 FILLER_0_33_139 ();
 FILLCELL_X1 FILLER_0_33_146 ();
 FILLCELL_X2 FILLER_0_33_150 ();
 FILLCELL_X2 FILLER_0_33_158 ();
 FILLCELL_X4 FILLER_0_33_173 ();
 FILLCELL_X1 FILLER_0_33_177 ();
 FILLCELL_X1 FILLER_0_33_216 ();
 FILLCELL_X8 FILLER_0_33_227 ();
 FILLCELL_X4 FILLER_0_33_247 ();
 FILLCELL_X8 FILLER_0_33_270 ();
 FILLCELL_X4 FILLER_0_33_278 ();
 FILLCELL_X2 FILLER_0_33_282 ();
 FILLCELL_X1 FILLER_0_33_284 ();
 FILLCELL_X1 FILLER_0_33_291 ();
 FILLCELL_X1 FILLER_0_33_296 ();
 FILLCELL_X1 FILLER_0_33_300 ();
 FILLCELL_X1 FILLER_0_33_305 ();
 FILLCELL_X2 FILLER_0_33_315 ();
 FILLCELL_X8 FILLER_0_33_326 ();
 FILLCELL_X4 FILLER_0_33_334 ();
 FILLCELL_X2 FILLER_0_33_338 ();
 FILLCELL_X1 FILLER_0_33_340 ();
 FILLCELL_X4 FILLER_0_33_351 ();
 FILLCELL_X1 FILLER_0_33_355 ();
 FILLCELL_X1 FILLER_0_33_367 ();
 FILLCELL_X4 FILLER_0_33_384 ();
 FILLCELL_X2 FILLER_0_34_1 ();
 FILLCELL_X1 FILLER_0_34_3 ();
 FILLCELL_X8 FILLER_0_34_7 ();
 FILLCELL_X4 FILLER_0_34_15 ();
 FILLCELL_X1 FILLER_0_34_19 ();
 FILLCELL_X1 FILLER_0_34_22 ();
 FILLCELL_X16 FILLER_0_34_32 ();
 FILLCELL_X2 FILLER_0_34_48 ();
 FILLCELL_X1 FILLER_0_34_50 ();
 FILLCELL_X1 FILLER_0_34_74 ();
 FILLCELL_X4 FILLER_0_34_104 ();
 FILLCELL_X2 FILLER_0_34_114 ();
 FILLCELL_X1 FILLER_0_34_116 ();
 FILLCELL_X1 FILLER_0_34_119 ();
 FILLCELL_X1 FILLER_0_34_129 ();
 FILLCELL_X2 FILLER_0_34_136 ();
 FILLCELL_X2 FILLER_0_34_148 ();
 FILLCELL_X1 FILLER_0_34_150 ();
 FILLCELL_X2 FILLER_0_34_163 ();
 FILLCELL_X1 FILLER_0_34_178 ();
 FILLCELL_X1 FILLER_0_34_187 ();
 FILLCELL_X1 FILLER_0_34_191 ();
 FILLCELL_X1 FILLER_0_34_198 ();
 FILLCELL_X2 FILLER_0_34_202 ();
 FILLCELL_X2 FILLER_0_34_208 ();
 FILLCELL_X1 FILLER_0_34_210 ();
 FILLCELL_X2 FILLER_0_34_224 ();
 FILLCELL_X1 FILLER_0_34_234 ();
 FILLCELL_X8 FILLER_0_34_245 ();
 FILLCELL_X4 FILLER_0_34_253 ();
 FILLCELL_X2 FILLER_0_34_257 ();
 FILLCELL_X2 FILLER_0_34_265 ();
 FILLCELL_X8 FILLER_0_34_271 ();
 FILLCELL_X2 FILLER_0_34_279 ();
 FILLCELL_X1 FILLER_0_34_281 ();
 FILLCELL_X1 FILLER_0_34_300 ();
 FILLCELL_X8 FILLER_0_34_304 ();
 FILLCELL_X2 FILLER_0_34_312 ();
 FILLCELL_X8 FILLER_0_34_333 ();
 FILLCELL_X16 FILLER_0_34_347 ();
 FILLCELL_X2 FILLER_0_34_363 ();
 FILLCELL_X1 FILLER_0_34_365 ();
 FILLCELL_X8 FILLER_0_34_379 ();
 FILLCELL_X1 FILLER_0_34_387 ();
 FILLCELL_X4 FILLER_0_35_1 ();
 FILLCELL_X1 FILLER_0_35_5 ();
 FILLCELL_X2 FILLER_0_35_9 ();
 FILLCELL_X1 FILLER_0_35_11 ();
 FILLCELL_X8 FILLER_0_35_37 ();
 FILLCELL_X2 FILLER_0_35_45 ();
 FILLCELL_X1 FILLER_0_35_55 ();
 FILLCELL_X1 FILLER_0_35_59 ();
 FILLCELL_X1 FILLER_0_35_69 ();
 FILLCELL_X1 FILLER_0_35_74 ();
 FILLCELL_X2 FILLER_0_35_81 ();
 FILLCELL_X1 FILLER_0_35_89 ();
 FILLCELL_X2 FILLER_0_35_94 ();
 FILLCELL_X2 FILLER_0_35_120 ();
 FILLCELL_X4 FILLER_0_35_132 ();
 FILLCELL_X1 FILLER_0_35_136 ();
 FILLCELL_X1 FILLER_0_35_160 ();
 FILLCELL_X1 FILLER_0_35_177 ();
 FILLCELL_X4 FILLER_0_35_189 ();
 FILLCELL_X8 FILLER_0_35_202 ();
 FILLCELL_X2 FILLER_0_35_210 ();
 FILLCELL_X1 FILLER_0_35_212 ();
 FILLCELL_X1 FILLER_0_35_243 ();
 FILLCELL_X2 FILLER_0_35_253 ();
 FILLCELL_X1 FILLER_0_35_255 ();
 FILLCELL_X2 FILLER_0_35_286 ();
 FILLCELL_X1 FILLER_0_35_288 ();
 FILLCELL_X4 FILLER_0_35_310 ();
 FILLCELL_X1 FILLER_0_35_325 ();
 FILLCELL_X4 FILLER_0_35_341 ();
 FILLCELL_X1 FILLER_0_35_351 ();
 FILLCELL_X1 FILLER_0_35_355 ();
 FILLCELL_X4 FILLER_0_35_378 ();
 FILLCELL_X2 FILLER_0_36_43 ();
 FILLCELL_X2 FILLER_0_36_57 ();
 FILLCELL_X4 FILLER_0_36_103 ();
 FILLCELL_X2 FILLER_0_36_107 ();
 FILLCELL_X1 FILLER_0_36_119 ();
 FILLCELL_X1 FILLER_0_36_123 ();
 FILLCELL_X1 FILLER_0_36_133 ();
 FILLCELL_X1 FILLER_0_36_151 ();
 FILLCELL_X2 FILLER_0_36_179 ();
 FILLCELL_X2 FILLER_0_36_201 ();
 FILLCELL_X4 FILLER_0_36_210 ();
 FILLCELL_X1 FILLER_0_36_214 ();
 FILLCELL_X4 FILLER_0_36_225 ();
 FILLCELL_X1 FILLER_0_36_233 ();
 FILLCELL_X2 FILLER_0_36_240 ();
 FILLCELL_X2 FILLER_0_36_246 ();
 FILLCELL_X2 FILLER_0_36_252 ();
 FILLCELL_X1 FILLER_0_36_254 ();
 FILLCELL_X1 FILLER_0_36_262 ();
 FILLCELL_X4 FILLER_0_36_284 ();
 FILLCELL_X1 FILLER_0_36_288 ();
 FILLCELL_X8 FILLER_0_36_301 ();
 FILLCELL_X4 FILLER_0_36_309 ();
 FILLCELL_X1 FILLER_0_36_313 ();
 FILLCELL_X1 FILLER_0_36_340 ();
 FILLCELL_X1 FILLER_0_36_345 ();
 FILLCELL_X1 FILLER_0_36_351 ();
 FILLCELL_X1 FILLER_0_36_358 ();
 FILLCELL_X1 FILLER_0_36_381 ();
 FILLCELL_X2 FILLER_0_37_28 ();
 FILLCELL_X1 FILLER_0_37_30 ();
 FILLCELL_X1 FILLER_0_37_34 ();
 FILLCELL_X2 FILLER_0_37_38 ();
 FILLCELL_X2 FILLER_0_37_44 ();
 FILLCELL_X1 FILLER_0_37_46 ();
 FILLCELL_X1 FILLER_0_37_59 ();
 FILLCELL_X1 FILLER_0_37_69 ();
 FILLCELL_X2 FILLER_0_37_85 ();
 FILLCELL_X2 FILLER_0_37_118 ();
 FILLCELL_X8 FILLER_0_37_126 ();
 FILLCELL_X4 FILLER_0_37_140 ();
 FILLCELL_X8 FILLER_0_37_148 ();
 FILLCELL_X4 FILLER_0_37_156 ();
 FILLCELL_X2 FILLER_0_37_160 ();
 FILLCELL_X1 FILLER_0_37_162 ();
 FILLCELL_X2 FILLER_0_37_176 ();
 FILLCELL_X4 FILLER_0_37_185 ();
 FILLCELL_X8 FILLER_0_37_199 ();
 FILLCELL_X4 FILLER_0_37_207 ();
 FILLCELL_X1 FILLER_0_37_211 ();
 FILLCELL_X8 FILLER_0_37_218 ();
 FILLCELL_X2 FILLER_0_37_226 ();
 FILLCELL_X2 FILLER_0_37_244 ();
 FILLCELL_X1 FILLER_0_37_260 ();
 FILLCELL_X4 FILLER_0_37_273 ();
 FILLCELL_X1 FILLER_0_37_277 ();
 FILLCELL_X2 FILLER_0_37_295 ();
 FILLCELL_X4 FILLER_0_37_313 ();
 FILLCELL_X1 FILLER_0_37_317 ();
 FILLCELL_X1 FILLER_0_37_326 ();
 FILLCELL_X1 FILLER_0_37_332 ();
 FILLCELL_X1 FILLER_0_37_339 ();
 FILLCELL_X1 FILLER_0_37_349 ();
 FILLCELL_X2 FILLER_0_37_353 ();
 FILLCELL_X1 FILLER_0_37_355 ();
 FILLCELL_X1 FILLER_0_37_357 ();
 FILLCELL_X1 FILLER_0_37_364 ();
 FILLCELL_X2 FILLER_0_37_371 ();
 FILLCELL_X4 FILLER_0_37_380 ();
 FILLCELL_X8 FILLER_0_38_1 ();
 FILLCELL_X4 FILLER_0_38_9 ();
 FILLCELL_X2 FILLER_0_38_25 ();
 FILLCELL_X1 FILLER_0_38_36 ();
 FILLCELL_X1 FILLER_0_38_41 ();
 FILLCELL_X1 FILLER_0_38_45 ();
 FILLCELL_X4 FILLER_0_38_55 ();
 FILLCELL_X2 FILLER_0_38_59 ();
 FILLCELL_X1 FILLER_0_38_83 ();
 FILLCELL_X1 FILLER_0_38_88 ();
 FILLCELL_X4 FILLER_0_38_90 ();
 FILLCELL_X1 FILLER_0_38_118 ();
 FILLCELL_X2 FILLER_0_38_125 ();
 FILLCELL_X2 FILLER_0_38_153 ();
 FILLCELL_X16 FILLER_0_38_158 ();
 FILLCELL_X4 FILLER_0_38_180 ();
 FILLCELL_X4 FILLER_0_38_187 ();
 FILLCELL_X1 FILLER_0_38_191 ();
 FILLCELL_X1 FILLER_0_38_198 ();
 FILLCELL_X2 FILLER_0_38_202 ();
 FILLCELL_X4 FILLER_0_38_210 ();
 FILLCELL_X2 FILLER_0_38_217 ();
 FILLCELL_X4 FILLER_0_38_225 ();
 FILLCELL_X1 FILLER_0_38_235 ();
 FILLCELL_X1 FILLER_0_38_247 ();
 FILLCELL_X2 FILLER_0_38_260 ();
 FILLCELL_X2 FILLER_0_38_268 ();
 FILLCELL_X1 FILLER_0_38_270 ();
 FILLCELL_X2 FILLER_0_38_277 ();
 FILLCELL_X1 FILLER_0_38_285 ();
 FILLCELL_X2 FILLER_0_38_289 ();
 FILLCELL_X4 FILLER_0_38_294 ();
 FILLCELL_X1 FILLER_0_38_298 ();
 FILLCELL_X2 FILLER_0_38_334 ();
 FILLCELL_X1 FILLER_0_38_336 ();
 FILLCELL_X2 FILLER_0_38_343 ();
 FILLCELL_X1 FILLER_0_38_377 ();
 FILLCELL_X4 FILLER_0_38_384 ();
 FILLCELL_X4 FILLER_0_39_1 ();
 FILLCELL_X2 FILLER_0_39_5 ();
 FILLCELL_X1 FILLER_0_39_7 ();
 FILLCELL_X2 FILLER_0_39_32 ();
 FILLCELL_X1 FILLER_0_39_51 ();
 FILLCELL_X4 FILLER_0_39_55 ();
 FILLCELL_X2 FILLER_0_39_59 ();
 FILLCELL_X2 FILLER_0_39_76 ();
 FILLCELL_X1 FILLER_0_39_78 ();
 FILLCELL_X4 FILLER_0_39_99 ();
 FILLCELL_X2 FILLER_0_39_103 ();
 FILLCELL_X1 FILLER_0_39_105 ();
 FILLCELL_X1 FILLER_0_39_128 ();
 FILLCELL_X4 FILLER_0_39_132 ();
 FILLCELL_X4 FILLER_0_39_159 ();
 FILLCELL_X2 FILLER_0_39_163 ();
 FILLCELL_X1 FILLER_0_39_165 ();
 FILLCELL_X2 FILLER_0_39_175 ();
 FILLCELL_X1 FILLER_0_39_177 ();
 FILLCELL_X4 FILLER_0_39_194 ();
 FILLCELL_X2 FILLER_0_39_211 ();
 FILLCELL_X2 FILLER_0_39_236 ();
 FILLCELL_X1 FILLER_0_39_260 ();
 FILLCELL_X1 FILLER_0_39_271 ();
 FILLCELL_X1 FILLER_0_39_284 ();
 FILLCELL_X1 FILLER_0_39_292 ();
 FILLCELL_X4 FILLER_0_39_320 ();
 FILLCELL_X4 FILLER_0_39_336 ();
 FILLCELL_X1 FILLER_0_39_355 ();
 FILLCELL_X1 FILLER_0_39_357 ();
 FILLCELL_X1 FILLER_0_39_361 ();
 FILLCELL_X1 FILLER_0_39_368 ();
 FILLCELL_X1 FILLER_0_39_371 ();
 FILLCELL_X2 FILLER_0_39_375 ();
 FILLCELL_X1 FILLER_0_39_377 ();
 FILLCELL_X4 FILLER_0_39_382 ();
 FILLCELL_X2 FILLER_0_39_386 ();
 FILLCELL_X4 FILLER_0_40_1 ();
 FILLCELL_X2 FILLER_0_40_5 ();
 FILLCELL_X4 FILLER_0_40_38 ();
 FILLCELL_X2 FILLER_0_40_42 ();
 FILLCELL_X1 FILLER_0_40_58 ();
 FILLCELL_X2 FILLER_0_40_93 ();
 FILLCELL_X1 FILLER_0_40_95 ();
 FILLCELL_X1 FILLER_0_40_105 ();
 FILLCELL_X1 FILLER_0_40_112 ();
 FILLCELL_X2 FILLER_0_40_117 ();
 FILLCELL_X4 FILLER_0_40_129 ();
 FILLCELL_X2 FILLER_0_40_133 ();
 FILLCELL_X1 FILLER_0_40_135 ();
 FILLCELL_X1 FILLER_0_40_146 ();
 FILLCELL_X4 FILLER_0_40_150 ();
 FILLCELL_X2 FILLER_0_40_154 ();
 FILLCELL_X1 FILLER_0_40_166 ();
 FILLCELL_X1 FILLER_0_40_173 ();
 FILLCELL_X2 FILLER_0_40_193 ();
 FILLCELL_X2 FILLER_0_40_207 ();
 FILLCELL_X1 FILLER_0_40_209 ();
 FILLCELL_X1 FILLER_0_40_225 ();
 FILLCELL_X1 FILLER_0_40_229 ();
 FILLCELL_X1 FILLER_0_40_234 ();
 FILLCELL_X1 FILLER_0_40_238 ();
 FILLCELL_X1 FILLER_0_40_243 ();
 FILLCELL_X4 FILLER_0_40_263 ();
 FILLCELL_X2 FILLER_0_40_268 ();
 FILLCELL_X8 FILLER_0_40_279 ();
 FILLCELL_X1 FILLER_0_40_287 ();
 FILLCELL_X1 FILLER_0_40_290 ();
 FILLCELL_X1 FILLER_0_40_297 ();
 FILLCELL_X1 FILLER_0_40_306 ();
 FILLCELL_X2 FILLER_0_40_317 ();
 FILLCELL_X1 FILLER_0_40_322 ();
 FILLCELL_X1 FILLER_0_40_330 ();
 FILLCELL_X1 FILLER_0_40_335 ();
 FILLCELL_X1 FILLER_0_40_345 ();
 FILLCELL_X2 FILLER_0_40_352 ();
 FILLCELL_X2 FILLER_0_40_364 ();
 FILLCELL_X1 FILLER_0_40_366 ();
 FILLCELL_X8 FILLER_0_40_376 ();
 FILLCELL_X4 FILLER_0_40_384 ();
 FILLCELL_X1 FILLER_0_41_1 ();
 FILLCELL_X1 FILLER_0_41_21 ();
 FILLCELL_X2 FILLER_0_41_53 ();
 FILLCELL_X1 FILLER_0_41_59 ();
 FILLCELL_X1 FILLER_0_41_63 ();
 FILLCELL_X1 FILLER_0_41_81 ();
 FILLCELL_X2 FILLER_0_41_86 ();
 FILLCELL_X2 FILLER_0_41_116 ();
 FILLCELL_X8 FILLER_0_41_127 ();
 FILLCELL_X1 FILLER_0_41_144 ();
 FILLCELL_X4 FILLER_0_41_150 ();
 FILLCELL_X1 FILLER_0_41_154 ();
 FILLCELL_X1 FILLER_0_41_161 ();
 FILLCELL_X2 FILLER_0_41_179 ();
 FILLCELL_X4 FILLER_0_41_193 ();
 FILLCELL_X1 FILLER_0_41_197 ();
 FILLCELL_X8 FILLER_0_41_204 ();
 FILLCELL_X4 FILLER_0_41_212 ();
 FILLCELL_X2 FILLER_0_41_216 ();
 FILLCELL_X1 FILLER_0_41_218 ();
 FILLCELL_X2 FILLER_0_41_232 ();
 FILLCELL_X1 FILLER_0_41_252 ();
 FILLCELL_X1 FILLER_0_41_256 ();
 FILLCELL_X1 FILLER_0_41_263 ();
 FILLCELL_X1 FILLER_0_41_268 ();
 FILLCELL_X1 FILLER_0_41_279 ();
 FILLCELL_X1 FILLER_0_41_292 ();
 FILLCELL_X2 FILLER_0_41_296 ();
 FILLCELL_X1 FILLER_0_41_298 ();
 FILLCELL_X1 FILLER_0_41_309 ();
 FILLCELL_X1 FILLER_0_41_313 ();
 FILLCELL_X1 FILLER_0_41_331 ();
 FILLCELL_X1 FILLER_0_41_341 ();
 FILLCELL_X1 FILLER_0_41_345 ();
 FILLCELL_X1 FILLER_0_41_352 ();
 FILLCELL_X1 FILLER_0_41_367 ();
 FILLCELL_X8 FILLER_0_41_374 ();
 FILLCELL_X4 FILLER_0_41_382 ();
 FILLCELL_X2 FILLER_0_41_386 ();
 FILLCELL_X4 FILLER_0_42_1 ();
 FILLCELL_X2 FILLER_0_42_37 ();
 FILLCELL_X1 FILLER_0_42_39 ();
 FILLCELL_X4 FILLER_0_42_52 ();
 FILLCELL_X1 FILLER_0_42_56 ();
 FILLCELL_X1 FILLER_0_42_81 ();
 FILLCELL_X2 FILLER_0_42_86 ();
 FILLCELL_X1 FILLER_0_42_88 ();
 FILLCELL_X1 FILLER_0_42_90 ();
 FILLCELL_X2 FILLER_0_42_97 ();
 FILLCELL_X4 FILLER_0_42_102 ();
 FILLCELL_X1 FILLER_0_42_106 ();
 FILLCELL_X2 FILLER_0_42_137 ();
 FILLCELL_X2 FILLER_0_42_156 ();
 FILLCELL_X2 FILLER_0_42_167 ();
 FILLCELL_X1 FILLER_0_42_169 ();
 FILLCELL_X2 FILLER_0_42_174 ();
 FILLCELL_X1 FILLER_0_42_176 ();
 FILLCELL_X1 FILLER_0_42_183 ();
 FILLCELL_X4 FILLER_0_42_189 ();
 FILLCELL_X8 FILLER_0_42_210 ();
 FILLCELL_X2 FILLER_0_42_218 ();
 FILLCELL_X1 FILLER_0_42_220 ();
 FILLCELL_X4 FILLER_0_42_239 ();
 FILLCELL_X1 FILLER_0_42_243 ();
 FILLCELL_X8 FILLER_0_42_258 ();
 FILLCELL_X1 FILLER_0_42_266 ();
 FILLCELL_X2 FILLER_0_42_268 ();
 FILLCELL_X1 FILLER_0_42_276 ();
 FILLCELL_X1 FILLER_0_42_281 ();
 FILLCELL_X4 FILLER_0_42_293 ();
 FILLCELL_X2 FILLER_0_42_309 ();
 FILLCELL_X2 FILLER_0_42_332 ();
 FILLCELL_X1 FILLER_0_42_337 ();
 FILLCELL_X4 FILLER_0_42_347 ();
 FILLCELL_X4 FILLER_0_42_354 ();
 FILLCELL_X2 FILLER_0_42_358 ();
 FILLCELL_X8 FILLER_0_42_373 ();
 FILLCELL_X4 FILLER_0_42_381 ();
 FILLCELL_X2 FILLER_0_42_385 ();
 FILLCELL_X1 FILLER_0_42_387 ();
 FILLCELL_X2 FILLER_0_43_1 ();
 FILLCELL_X1 FILLER_0_43_3 ();
 FILLCELL_X1 FILLER_0_43_11 ();
 FILLCELL_X1 FILLER_0_43_15 ();
 FILLCELL_X1 FILLER_0_43_20 ();
 FILLCELL_X2 FILLER_0_43_33 ();
 FILLCELL_X1 FILLER_0_43_39 ();
 FILLCELL_X1 FILLER_0_43_46 ();
 FILLCELL_X2 FILLER_0_43_51 ();
 FILLCELL_X1 FILLER_0_43_53 ();
 FILLCELL_X4 FILLER_0_43_57 ();
 FILLCELL_X2 FILLER_0_43_61 ();
 FILLCELL_X2 FILLER_0_43_111 ();
 FILLCELL_X1 FILLER_0_43_129 ();
 FILLCELL_X1 FILLER_0_43_136 ();
 FILLCELL_X1 FILLER_0_43_144 ();
 FILLCELL_X8 FILLER_0_43_147 ();
 FILLCELL_X4 FILLER_0_43_155 ();
 FILLCELL_X1 FILLER_0_43_159 ();
 FILLCELL_X4 FILLER_0_43_166 ();
 FILLCELL_X1 FILLER_0_43_170 ();
 FILLCELL_X8 FILLER_0_43_185 ();
 FILLCELL_X8 FILLER_0_43_196 ();
 FILLCELL_X4 FILLER_0_43_221 ();
 FILLCELL_X2 FILLER_0_43_225 ();
 FILLCELL_X2 FILLER_0_43_233 ();
 FILLCELL_X1 FILLER_0_43_243 ();
 FILLCELL_X1 FILLER_0_43_248 ();
 FILLCELL_X2 FILLER_0_43_253 ();
 FILLCELL_X1 FILLER_0_43_255 ();
 FILLCELL_X1 FILLER_0_43_273 ();
 FILLCELL_X1 FILLER_0_43_296 ();
 FILLCELL_X1 FILLER_0_43_300 ();
 FILLCELL_X1 FILLER_0_43_305 ();
 FILLCELL_X1 FILLER_0_43_309 ();
 FILLCELL_X1 FILLER_0_43_330 ();
 FILLCELL_X16 FILLER_0_43_339 ();
 FILLCELL_X1 FILLER_0_43_355 ();
 FILLCELL_X2 FILLER_0_43_386 ();
 FILLCELL_X1 FILLER_0_44_18 ();
 FILLCELL_X2 FILLER_0_44_24 ();
 FILLCELL_X2 FILLER_0_44_35 ();
 FILLCELL_X2 FILLER_0_44_43 ();
 FILLCELL_X1 FILLER_0_44_45 ();
 FILLCELL_X2 FILLER_0_44_52 ();
 FILLCELL_X1 FILLER_0_44_54 ();
 FILLCELL_X2 FILLER_0_44_61 ();
 FILLCELL_X4 FILLER_0_44_73 ();
 FILLCELL_X1 FILLER_0_44_77 ();
 FILLCELL_X4 FILLER_0_44_82 ();
 FILLCELL_X1 FILLER_0_44_103 ();
 FILLCELL_X2 FILLER_0_44_110 ();
 FILLCELL_X1 FILLER_0_44_112 ();
 FILLCELL_X2 FILLER_0_44_119 ();
 FILLCELL_X2 FILLER_0_44_130 ();
 FILLCELL_X1 FILLER_0_44_132 ();
 FILLCELL_X2 FILLER_0_44_155 ();
 FILLCELL_X2 FILLER_0_44_172 ();
 FILLCELL_X1 FILLER_0_44_174 ();
 FILLCELL_X2 FILLER_0_44_206 ();
 FILLCELL_X8 FILLER_0_44_216 ();
 FILLCELL_X4 FILLER_0_44_224 ();
 FILLCELL_X1 FILLER_0_44_249 ();
 FILLCELL_X4 FILLER_0_44_268 ();
 FILLCELL_X2 FILLER_0_44_272 ();
 FILLCELL_X1 FILLER_0_44_326 ();
 FILLCELL_X1 FILLER_0_44_331 ();
 FILLCELL_X1 FILLER_0_44_337 ();
 FILLCELL_X8 FILLER_0_44_355 ();
 FILLCELL_X4 FILLER_0_44_363 ();
 FILLCELL_X2 FILLER_0_44_367 ();
 FILLCELL_X8 FILLER_0_44_375 ();
 FILLCELL_X4 FILLER_0_44_383 ();
 FILLCELL_X1 FILLER_0_44_387 ();
 FILLCELL_X8 FILLER_0_45_1 ();
 FILLCELL_X2 FILLER_0_45_9 ();
 FILLCELL_X1 FILLER_0_45_26 ();
 FILLCELL_X1 FILLER_0_45_30 ();
 FILLCELL_X1 FILLER_0_45_34 ();
 FILLCELL_X1 FILLER_0_45_42 ();
 FILLCELL_X8 FILLER_0_45_53 ();
 FILLCELL_X2 FILLER_0_45_61 ();
 FILLCELL_X1 FILLER_0_45_78 ();
 FILLCELL_X1 FILLER_0_45_96 ();
 FILLCELL_X2 FILLER_0_45_101 ();
 FILLCELL_X1 FILLER_0_45_103 ();
 FILLCELL_X1 FILLER_0_45_127 ();
 FILLCELL_X4 FILLER_0_45_132 ();
 FILLCELL_X1 FILLER_0_45_136 ();
 FILLCELL_X8 FILLER_0_45_143 ();
 FILLCELL_X1 FILLER_0_45_151 ();
 FILLCELL_X1 FILLER_0_45_160 ();
 FILLCELL_X1 FILLER_0_45_164 ();
 FILLCELL_X1 FILLER_0_45_173 ();
 FILLCELL_X2 FILLER_0_45_179 ();
 FILLCELL_X1 FILLER_0_45_185 ();
 FILLCELL_X2 FILLER_0_45_211 ();
 FILLCELL_X1 FILLER_0_45_216 ();
 FILLCELL_X4 FILLER_0_45_220 ();
 FILLCELL_X1 FILLER_0_45_232 ();
 FILLCELL_X1 FILLER_0_45_267 ();
 FILLCELL_X2 FILLER_0_45_277 ();
 FILLCELL_X1 FILLER_0_45_279 ();
 FILLCELL_X1 FILLER_0_45_292 ();
 FILLCELL_X1 FILLER_0_45_352 ();
 FILLCELL_X16 FILLER_0_45_361 ();
 FILLCELL_X8 FILLER_0_45_377 ();
 FILLCELL_X2 FILLER_0_45_385 ();
 FILLCELL_X1 FILLER_0_45_387 ();
 FILLCELL_X8 FILLER_0_46_1 ();
 FILLCELL_X4 FILLER_0_46_9 ();
 FILLCELL_X1 FILLER_0_46_13 ();
 FILLCELL_X2 FILLER_0_46_27 ();
 FILLCELL_X1 FILLER_0_46_33 ();
 FILLCELL_X1 FILLER_0_46_42 ();
 FILLCELL_X1 FILLER_0_46_49 ();
 FILLCELL_X2 FILLER_0_46_56 ();
 FILLCELL_X2 FILLER_0_46_64 ();
 FILLCELL_X1 FILLER_0_46_68 ();
 FILLCELL_X1 FILLER_0_46_74 ();
 FILLCELL_X1 FILLER_0_46_82 ();
 FILLCELL_X4 FILLER_0_46_94 ();
 FILLCELL_X1 FILLER_0_46_98 ();
 FILLCELL_X2 FILLER_0_46_105 ();
 FILLCELL_X1 FILLER_0_46_107 ();
 FILLCELL_X2 FILLER_0_46_122 ();
 FILLCELL_X1 FILLER_0_46_128 ();
 FILLCELL_X1 FILLER_0_46_134 ();
 FILLCELL_X1 FILLER_0_46_145 ();
 FILLCELL_X1 FILLER_0_46_154 ();
 FILLCELL_X1 FILLER_0_46_187 ();
 FILLCELL_X2 FILLER_0_46_202 ();
 FILLCELL_X1 FILLER_0_46_214 ();
 FILLCELL_X1 FILLER_0_46_261 ();
 FILLCELL_X1 FILLER_0_46_266 ();
 FILLCELL_X8 FILLER_0_46_273 ();
 FILLCELL_X4 FILLER_0_46_281 ();
 FILLCELL_X2 FILLER_0_46_285 ();
 FILLCELL_X4 FILLER_0_46_293 ();
 FILLCELL_X8 FILLER_0_46_303 ();
 FILLCELL_X1 FILLER_0_46_311 ();
 FILLCELL_X2 FILLER_0_46_330 ();
 FILLCELL_X2 FILLER_0_46_353 ();
 FILLCELL_X1 FILLER_0_46_355 ();
 FILLCELL_X16 FILLER_0_46_362 ();
 FILLCELL_X8 FILLER_0_46_378 ();
 FILLCELL_X2 FILLER_0_46_386 ();
 FILLCELL_X8 FILLER_0_47_1 ();
 FILLCELL_X4 FILLER_0_47_9 ();
 FILLCELL_X2 FILLER_0_47_13 ();
 FILLCELL_X1 FILLER_0_47_15 ();
 FILLCELL_X1 FILLER_0_47_19 ();
 FILLCELL_X4 FILLER_0_47_23 ();
 FILLCELL_X4 FILLER_0_47_39 ();
 FILLCELL_X2 FILLER_0_47_43 ();
 FILLCELL_X4 FILLER_0_47_58 ();
 FILLCELL_X2 FILLER_0_47_62 ();
 FILLCELL_X4 FILLER_0_47_103 ();
 FILLCELL_X4 FILLER_0_47_122 ();
 FILLCELL_X1 FILLER_0_47_126 ();
 FILLCELL_X2 FILLER_0_47_146 ();
 FILLCELL_X2 FILLER_0_47_158 ();
 FILLCELL_X2 FILLER_0_47_185 ();
 FILLCELL_X1 FILLER_0_47_187 ();
 FILLCELL_X1 FILLER_0_47_197 ();
 FILLCELL_X1 FILLER_0_47_216 ();
 FILLCELL_X1 FILLER_0_47_221 ();
 FILLCELL_X1 FILLER_0_47_226 ();
 FILLCELL_X1 FILLER_0_47_233 ();
 FILLCELL_X8 FILLER_0_47_236 ();
 FILLCELL_X4 FILLER_0_47_244 ();
 FILLCELL_X2 FILLER_0_47_248 ();
 FILLCELL_X8 FILLER_0_47_260 ();
 FILLCELL_X2 FILLER_0_47_268 ();
 FILLCELL_X2 FILLER_0_47_295 ();
 FILLCELL_X4 FILLER_0_47_303 ();
 FILLCELL_X2 FILLER_0_47_307 ();
 FILLCELL_X8 FILLER_0_47_313 ();
 FILLCELL_X1 FILLER_0_47_321 ();
 FILLCELL_X1 FILLER_0_47_332 ();
 FILLCELL_X1 FILLER_0_47_350 ();
 FILLCELL_X2 FILLER_0_47_354 ();
 FILLCELL_X16 FILLER_0_47_357 ();
 FILLCELL_X8 FILLER_0_47_373 ();
 FILLCELL_X4 FILLER_0_47_381 ();
 FILLCELL_X2 FILLER_0_47_385 ();
 FILLCELL_X1 FILLER_0_47_387 ();
 FILLCELL_X16 FILLER_0_48_1 ();
 FILLCELL_X1 FILLER_0_48_38 ();
 FILLCELL_X1 FILLER_0_48_47 ();
 FILLCELL_X1 FILLER_0_48_60 ();
 FILLCELL_X1 FILLER_0_48_65 ();
 FILLCELL_X1 FILLER_0_48_84 ();
 FILLCELL_X1 FILLER_0_48_88 ();
 FILLCELL_X4 FILLER_0_48_93 ();
 FILLCELL_X2 FILLER_0_48_97 ();
 FILLCELL_X1 FILLER_0_48_105 ();
 FILLCELL_X2 FILLER_0_48_112 ();
 FILLCELL_X1 FILLER_0_48_114 ();
 FILLCELL_X2 FILLER_0_48_130 ();
 FILLCELL_X8 FILLER_0_48_144 ();
 FILLCELL_X1 FILLER_0_48_158 ();
 FILLCELL_X2 FILLER_0_48_165 ();
 FILLCELL_X1 FILLER_0_48_169 ();
 FILLCELL_X2 FILLER_0_48_173 ();
 FILLCELL_X1 FILLER_0_48_181 ();
 FILLCELL_X8 FILLER_0_48_215 ();
 FILLCELL_X2 FILLER_0_48_223 ();
 FILLCELL_X1 FILLER_0_48_225 ();
 FILLCELL_X2 FILLER_0_48_249 ();
 FILLCELL_X1 FILLER_0_48_255 ();
 FILLCELL_X2 FILLER_0_48_265 ();
 FILLCELL_X4 FILLER_0_48_274 ();
 FILLCELL_X2 FILLER_0_48_278 ();
 FILLCELL_X1 FILLER_0_48_280 ();
 FILLCELL_X1 FILLER_0_48_286 ();
 FILLCELL_X1 FILLER_0_48_299 ();
 FILLCELL_X2 FILLER_0_48_305 ();
 FILLCELL_X1 FILLER_0_48_307 ();
 FILLCELL_X1 FILLER_0_48_314 ();
 FILLCELL_X1 FILLER_0_48_318 ();
 FILLCELL_X1 FILLER_0_48_322 ();
 FILLCELL_X2 FILLER_0_48_329 ();
 FILLCELL_X1 FILLER_0_48_331 ();
 FILLCELL_X2 FILLER_0_48_338 ();
 FILLCELL_X1 FILLER_0_48_346 ();
 FILLCELL_X32 FILLER_0_48_349 ();
 FILLCELL_X4 FILLER_0_48_381 ();
 FILLCELL_X2 FILLER_0_48_385 ();
 FILLCELL_X1 FILLER_0_48_387 ();
 FILLCELL_X16 FILLER_0_49_1 ();
 FILLCELL_X8 FILLER_0_49_17 ();
 FILLCELL_X2 FILLER_0_49_25 ();
 FILLCELL_X1 FILLER_0_49_27 ();
 FILLCELL_X1 FILLER_0_49_40 ();
 FILLCELL_X1 FILLER_0_49_49 ();
 FILLCELL_X2 FILLER_0_49_81 ();
 FILLCELL_X2 FILLER_0_49_93 ();
 FILLCELL_X1 FILLER_0_49_104 ();
 FILLCELL_X4 FILLER_0_49_111 ();
 FILLCELL_X2 FILLER_0_49_115 ();
 FILLCELL_X8 FILLER_0_49_122 ();
 FILLCELL_X2 FILLER_0_49_130 ();
 FILLCELL_X1 FILLER_0_49_132 ();
 FILLCELL_X4 FILLER_0_49_172 ();
 FILLCELL_X2 FILLER_0_49_176 ();
 FILLCELL_X1 FILLER_0_49_187 ();
 FILLCELL_X4 FILLER_0_49_191 ();
 FILLCELL_X1 FILLER_0_49_195 ();
 FILLCELL_X2 FILLER_0_49_222 ();
 FILLCELL_X1 FILLER_0_49_230 ();
 FILLCELL_X1 FILLER_0_49_244 ();
 FILLCELL_X4 FILLER_0_49_276 ();
 FILLCELL_X2 FILLER_0_49_280 ();
 FILLCELL_X1 FILLER_0_49_288 ();
 FILLCELL_X1 FILLER_0_49_294 ();
 FILLCELL_X1 FILLER_0_49_301 ();
 FILLCELL_X2 FILLER_0_49_308 ();
 FILLCELL_X16 FILLER_0_49_332 ();
 FILLCELL_X8 FILLER_0_49_348 ();
 FILLCELL_X16 FILLER_0_49_357 ();
 FILLCELL_X8 FILLER_0_49_373 ();
 FILLCELL_X4 FILLER_0_49_381 ();
 FILLCELL_X2 FILLER_0_49_385 ();
 FILLCELL_X1 FILLER_0_49_387 ();
 FILLCELL_X16 FILLER_0_50_1 ();
 FILLCELL_X8 FILLER_0_50_17 ();
 FILLCELL_X1 FILLER_0_50_25 ();
 FILLCELL_X2 FILLER_0_50_30 ();
 FILLCELL_X2 FILLER_0_50_47 ();
 FILLCELL_X2 FILLER_0_50_53 ();
 FILLCELL_X1 FILLER_0_50_55 ();
 FILLCELL_X2 FILLER_0_50_73 ();
 FILLCELL_X1 FILLER_0_50_75 ();
 FILLCELL_X2 FILLER_0_50_80 ();
 FILLCELL_X1 FILLER_0_50_82 ();
 FILLCELL_X2 FILLER_0_50_94 ();
 FILLCELL_X1 FILLER_0_50_111 ();
 FILLCELL_X1 FILLER_0_50_118 ();
 FILLCELL_X1 FILLER_0_50_125 ();
 FILLCELL_X1 FILLER_0_50_132 ();
 FILLCELL_X2 FILLER_0_50_135 ();
 FILLCELL_X1 FILLER_0_50_157 ();
 FILLCELL_X8 FILLER_0_50_167 ();
 FILLCELL_X4 FILLER_0_50_175 ();
 FILLCELL_X2 FILLER_0_50_179 ();
 FILLCELL_X1 FILLER_0_50_181 ();
 FILLCELL_X4 FILLER_0_50_205 ();
 FILLCELL_X1 FILLER_0_50_209 ();
 FILLCELL_X1 FILLER_0_50_216 ();
 FILLCELL_X1 FILLER_0_50_223 ();
 FILLCELL_X1 FILLER_0_50_227 ();
 FILLCELL_X1 FILLER_0_50_232 ();
 FILLCELL_X1 FILLER_0_50_236 ();
 FILLCELL_X1 FILLER_0_50_243 ();
 FILLCELL_X2 FILLER_0_50_257 ();
 FILLCELL_X1 FILLER_0_50_262 ();
 FILLCELL_X1 FILLER_0_50_268 ();
 FILLCELL_X2 FILLER_0_50_275 ();
 FILLCELL_X2 FILLER_0_50_292 ();
 FILLCELL_X4 FILLER_0_50_298 ();
 FILLCELL_X2 FILLER_0_50_302 ();
 FILLCELL_X1 FILLER_0_50_304 ();
 FILLCELL_X32 FILLER_0_50_331 ();
 FILLCELL_X8 FILLER_0_50_363 ();
 FILLCELL_X8 FILLER_0_50_375 ();
 FILLCELL_X4 FILLER_0_50_383 ();
 FILLCELL_X1 FILLER_0_50_387 ();
 FILLCELL_X32 FILLER_0_51_1 ();
 FILLCELL_X16 FILLER_0_51_50 ();
 FILLCELL_X4 FILLER_0_51_66 ();
 FILLCELL_X2 FILLER_0_51_70 ();
 FILLCELL_X1 FILLER_0_51_88 ();
 FILLCELL_X1 FILLER_0_51_90 ();
 FILLCELL_X1 FILLER_0_51_115 ();
 FILLCELL_X2 FILLER_0_51_118 ();
 FILLCELL_X1 FILLER_0_51_124 ();
 FILLCELL_X4 FILLER_0_51_128 ();
 FILLCELL_X2 FILLER_0_51_132 ();
 FILLCELL_X1 FILLER_0_51_141 ();
 FILLCELL_X4 FILLER_0_51_149 ();
 FILLCELL_X1 FILLER_0_51_177 ();
 FILLCELL_X1 FILLER_0_51_179 ();
 FILLCELL_X1 FILLER_0_51_183 ();
 FILLCELL_X16 FILLER_0_51_187 ();
 FILLCELL_X8 FILLER_0_51_203 ();
 FILLCELL_X4 FILLER_0_51_211 ();
 FILLCELL_X2 FILLER_0_51_215 ();
 FILLCELL_X1 FILLER_0_51_221 ();
 FILLCELL_X1 FILLER_0_51_228 ();
 FILLCELL_X1 FILLER_0_51_232 ();
 FILLCELL_X1 FILLER_0_51_239 ();
 FILLCELL_X8 FILLER_0_51_253 ();
 FILLCELL_X2 FILLER_0_51_286 ();
 FILLCELL_X16 FILLER_0_51_297 ();
 FILLCELL_X4 FILLER_0_51_313 ();
 FILLCELL_X16 FILLER_0_51_332 ();
 FILLCELL_X8 FILLER_0_51_348 ();
 FILLCELL_X16 FILLER_0_51_357 ();
 FILLCELL_X8 FILLER_0_51_373 ();
 FILLCELL_X4 FILLER_0_51_381 ();
 FILLCELL_X2 FILLER_0_51_385 ();
 FILLCELL_X1 FILLER_0_51_387 ();
endmodule
