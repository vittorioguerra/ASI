module enfasi (clk,
    rst,
    q,
    z);
 input clk;
 input rst;
 output [11:0] q;
 input [10:0] z;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire \aso.p[0] ;
 wire \aso.p[10] ;
 wire \aso.p[11] ;
 wire \aso.p[1] ;
 wire \aso.p[2] ;
 wire \aso.p[3] ;
 wire \aso.p[4] ;
 wire \aso.p[5] ;
 wire \aso.p[6] ;
 wire \aso.p[7] ;
 wire \aso.p[8] ;
 wire \aso.p[9] ;
 wire \aso.z0[0] ;
 wire \aso.z0[10] ;
 wire \aso.z0[1] ;
 wire \aso.z0[2] ;
 wire \aso.z0[3] ;
 wire \aso.z0[4] ;
 wire \aso.z0[5] ;
 wire \aso.z0[6] ;
 wire \aso.z0[7] ;
 wire \aso.z0[8] ;
 wire \aso.z0[9] ;
 wire \aso.z1[0] ;
 wire \aso.z1[10] ;
 wire \aso.z1[1] ;
 wire \aso.z1[2] ;
 wire \aso.z1[3] ;
 wire \aso.z1[4] ;
 wire \aso.z1[5] ;
 wire \aso.z1[6] ;
 wire \aso.z1[7] ;
 wire \aso.z1[8] ;
 wire \aso.z1[9] ;
 wire \aso.z2[0] ;
 wire \aso.z2[10] ;
 wire \aso.z2[1] ;
 wire \aso.z2[2] ;
 wire \aso.z2[3] ;
 wire \aso.z2[4] ;
 wire \aso.z2[5] ;
 wire \aso.z2[6] ;
 wire \aso.z2[7] ;
 wire \aso.z2[8] ;
 wire \aso.z2[9] ;
 wire \aso.z3[0] ;
 wire \aso.z3[10] ;
 wire \aso.z3[1] ;
 wire \aso.z3[2] ;
 wire \aso.z3[3] ;
 wire \aso.z3[4] ;
 wire \aso.z3[5] ;
 wire \aso.z3[6] ;
 wire \aso.z3[7] ;
 wire \aso.z3[8] ;
 wire \aso.z3[9] ;
 wire \aso.z4[0] ;
 wire \aso.z4[10] ;
 wire \aso.z4[1] ;
 wire \aso.z4[2] ;
 wire \aso.z4[3] ;
 wire \aso.z4[4] ;
 wire \aso.z4[5] ;
 wire \aso.z4[6] ;
 wire \aso.z4[7] ;
 wire \aso.z4[8] ;
 wire \aso.z4[9] ;
 wire \fir.p0[0] ;
 wire \fir.p0[10] ;
 wire \fir.p0[11] ;
 wire \fir.p0[1] ;
 wire \fir.p0[2] ;
 wire \fir.p0[3] ;
 wire \fir.p0[4] ;
 wire \fir.p0[5] ;
 wire \fir.p0[6] ;
 wire \fir.p0[7] ;
 wire \fir.p0[8] ;
 wire \fir.p0[9] ;
 wire \fir.p1[0] ;
 wire \fir.p1[10] ;
 wire \fir.p1[11] ;
 wire \fir.p1[1] ;
 wire \fir.p1[2] ;
 wire \fir.p1[3] ;
 wire \fir.p1[4] ;
 wire \fir.p1[5] ;
 wire \fir.p1[6] ;
 wire \fir.p1[7] ;
 wire \fir.p1[8] ;
 wire \fir.p1[9] ;
 wire \fir.p2[0] ;
 wire \fir.p2[10] ;
 wire \fir.p2[11] ;
 wire \fir.p2[1] ;
 wire \fir.p2[2] ;
 wire \fir.p2[3] ;
 wire \fir.p2[4] ;
 wire \fir.p2[5] ;
 wire \fir.p2[6] ;
 wire \fir.p2[7] ;
 wire \fir.p2[8] ;
 wire \fir.p2[9] ;
 wire \fir.p3[0] ;
 wire \fir.p3[10] ;
 wire \fir.p3[11] ;
 wire \fir.p3[1] ;
 wire \fir.p3[2] ;
 wire \fir.p3[3] ;
 wire \fir.p3[4] ;
 wire \fir.p3[5] ;
 wire \fir.p3[6] ;
 wire \fir.p3[7] ;
 wire \fir.p3[8] ;
 wire \fir.p3[9] ;
 wire \fir.p4[0] ;
 wire \fir.p4[10] ;
 wire \fir.p4[11] ;
 wire \fir.p4[1] ;
 wire \fir.p4[2] ;
 wire \fir.p4[3] ;
 wire \fir.p4[4] ;
 wire \fir.p4[5] ;
 wire \fir.p4[6] ;
 wire \fir.p4[7] ;
 wire \fir.p4[8] ;
 wire \fir.p4[9] ;
 wire \fir.p5[0] ;
 wire \fir.p5[10] ;
 wire \fir.p5[11] ;
 wire \fir.p5[1] ;
 wire \fir.p5[2] ;
 wire \fir.p5[3] ;
 wire \fir.p5[4] ;
 wire \fir.p5[5] ;
 wire \fir.p5[6] ;
 wire \fir.p5[7] ;
 wire \fir.p5[8] ;
 wire \fir.p5[9] ;
 wire \fir.p6[0] ;
 wire \fir.p6[10] ;
 wire \fir.p6[11] ;
 wire \fir.p6[1] ;
 wire \fir.p6[2] ;
 wire \fir.p6[3] ;
 wire \fir.p6[4] ;
 wire \fir.p6[5] ;
 wire \fir.p6[6] ;
 wire \fir.p6[7] ;
 wire \fir.p6[8] ;
 wire \fir.p6[9] ;
 wire \fir.p7[0] ;
 wire \fir.p7[10] ;
 wire \fir.p7[11] ;
 wire \fir.p7[1] ;
 wire \fir.p7[2] ;
 wire \fir.p7[3] ;
 wire \fir.p7[4] ;
 wire \fir.p7[5] ;
 wire \fir.p7[6] ;
 wire \fir.p7[7] ;
 wire \fir.p7[8] ;
 wire \fir.p7[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;

 INV_X1 _3802_ (.A(rst),
    .ZN(_2962_));
 NAND2_X1 _3803_ (.A1(\fir.p7[11] ),
    .A2(\fir.p7[9] ),
    .ZN(_2973_));
 NOR3_X1 _3804_ (.A1(_0037_),
    .A2(_0031_),
    .A3(_2973_),
    .ZN(_2984_));
 NAND2_X1 _3805_ (.A1(\fir.p1[0] ),
    .A2(\fir.p0[0] ),
    .ZN(_2995_));
 OR2_X1 _3806_ (.A1(\fir.p1[1] ),
    .A2(\fir.p1[0] ),
    .ZN(_3006_));
 NAND2_X1 _3807_ (.A1(\fir.p1[1] ),
    .A2(\fir.p1[0] ),
    .ZN(_3015_));
 NAND2_X1 _3808_ (.A1(_3006_),
    .A2(_3015_),
    .ZN(_3021_));
 XOR2_X1 _3809_ (.A(\fir.p0[1] ),
    .B(_3021_),
    .Z(_3030_));
 XOR2_X1 _3810_ (.A(_2995_),
    .B(_3030_),
    .Z(_3041_));
 NAND2_X1 _3811_ (.A1(\fir.p2[0] ),
    .A2(_3041_),
    .ZN(_3052_));
 NOR2_X1 _3812_ (.A1(_2995_),
    .A2(_3030_),
    .ZN(_3063_));
 NAND3_X1 _3813_ (.A1(\fir.p0[1] ),
    .A2(_3006_),
    .A3(_3015_),
    .ZN(_3069_));
 XOR2_X1 _3814_ (.A(\fir.p0[2] ),
    .B(\fir.p0[0] ),
    .Z(_3070_));
 XOR2_X1 _3815_ (.A(\fir.p1[2] ),
    .B(\fir.p1[1] ),
    .Z(_3071_));
 XNOR2_X1 _3816_ (.A(_3015_),
    .B(_3071_),
    .ZN(_3072_));
 XNOR2_X1 _3817_ (.A(_3070_),
    .B(_3072_),
    .ZN(_3073_));
 XNOR2_X1 _3818_ (.A(_3069_),
    .B(_3073_),
    .ZN(_3074_));
 XNOR2_X1 _3819_ (.A(_3063_),
    .B(_3074_),
    .ZN(_3075_));
 XNOR2_X1 _3820_ (.A(\fir.p2[1] ),
    .B(_3075_),
    .ZN(_3076_));
 NOR2_X1 _3821_ (.A1(_3052_),
    .A2(_3076_),
    .ZN(_3077_));
 NAND2_X1 _3822_ (.A1(\fir.p2[1] ),
    .A2(_3075_),
    .ZN(_3078_));
 NAND2_X1 _3823_ (.A1(_3070_),
    .A2(_3072_),
    .ZN(_3079_));
 NAND2_X1 _3824_ (.A1(\fir.p0[2] ),
    .A2(\fir.p0[0] ),
    .ZN(_3080_));
 XOR2_X1 _3825_ (.A(\fir.p0[3] ),
    .B(\fir.p0[1] ),
    .Z(_3081_));
 XNOR2_X1 _3826_ (.A(_3080_),
    .B(_3081_),
    .ZN(_3082_));
 NAND2_X1 _3827_ (.A1(\fir.p1[2] ),
    .A2(\fir.p1[1] ),
    .ZN(_3083_));
 XOR2_X1 _3828_ (.A(\fir.p1[3] ),
    .B(\fir.p1[2] ),
    .Z(_3084_));
 XNOR2_X1 _3829_ (.A(_3083_),
    .B(_3084_),
    .ZN(_3085_));
 XNOR2_X1 _3830_ (.A(_3082_),
    .B(_3085_),
    .ZN(_3086_));
 XNOR2_X1 _3831_ (.A(_3079_),
    .B(_3086_),
    .ZN(_3087_));
 OR3_X1 _3832_ (.A1(\fir.p1[2] ),
    .A2(_3015_),
    .A3(_3087_),
    .ZN(_3088_));
 OAI21_X1 _3833_ (.A(_3087_),
    .B1(_3015_),
    .B2(\fir.p1[2] ),
    .ZN(_3089_));
 AND2_X1 _3834_ (.A1(_3088_),
    .A2(_3089_),
    .ZN(_3090_));
 NOR2_X1 _3835_ (.A1(_3069_),
    .A2(_3073_),
    .ZN(_3091_));
 NOR3_X1 _3836_ (.A1(_2995_),
    .A2(_3030_),
    .A3(_3074_),
    .ZN(_3092_));
 NOR2_X1 _3837_ (.A1(_3091_),
    .A2(_3092_),
    .ZN(_3093_));
 XNOR2_X1 _3838_ (.A(_3090_),
    .B(_3093_),
    .ZN(_3094_));
 XOR2_X1 _3839_ (.A(\fir.p2[0] ),
    .B(_3094_),
    .Z(_3095_));
 NAND2_X1 _3840_ (.A1(\fir.p2[2] ),
    .A2(_3095_),
    .ZN(_3096_));
 INV_X1 _3841_ (.A(_3096_),
    .ZN(_3097_));
 NOR2_X1 _3842_ (.A1(\fir.p2[2] ),
    .A2(_3095_),
    .ZN(_3098_));
 OR2_X1 _3843_ (.A1(_3097_),
    .A2(_3098_),
    .ZN(_3099_));
 XOR2_X1 _3844_ (.A(_3078_),
    .B(_3099_),
    .Z(_3100_));
 XOR2_X1 _3845_ (.A(_3077_),
    .B(_3100_),
    .Z(_3101_));
 NAND2_X1 _3846_ (.A1(\fir.p4[3] ),
    .A2(_3101_),
    .ZN(_3102_));
 NAND2_X1 _3847_ (.A1(\fir.p2[0] ),
    .A2(_3094_),
    .ZN(_3103_));
 NAND2_X1 _3848_ (.A1(_3092_),
    .A2(_3090_),
    .ZN(_3104_));
 NAND2_X1 _3849_ (.A1(_3091_),
    .A2(_3090_),
    .ZN(_3105_));
 OAI21_X1 _3850_ (.A(_3088_),
    .B1(_3086_),
    .B2(_3079_),
    .ZN(_3106_));
 OR2_X1 _3851_ (.A1(\fir.p1[3] ),
    .A2(_3083_),
    .ZN(_3107_));
 NAND2_X1 _3852_ (.A1(_3082_),
    .A2(_3085_),
    .ZN(_3108_));
 AND3_X1 _3853_ (.A1(\fir.p0[2] ),
    .A2(\fir.p0[0] ),
    .A3(_3081_),
    .ZN(_3109_));
 NAND2_X1 _3854_ (.A1(\fir.p0[3] ),
    .A2(\fir.p0[1] ),
    .ZN(_3110_));
 XOR2_X1 _3855_ (.A(\fir.p0[4] ),
    .B(\fir.p0[2] ),
    .Z(_3111_));
 XNOR2_X1 _3856_ (.A(_3110_),
    .B(_3111_),
    .ZN(_3112_));
 XNOR2_X1 _3857_ (.A(\fir.p0[0] ),
    .B(_3112_),
    .ZN(_3113_));
 XNOR2_X1 _3858_ (.A(_3109_),
    .B(_3113_),
    .ZN(_3114_));
 NAND2_X1 _3859_ (.A1(\fir.p1[3] ),
    .A2(\fir.p1[2] ),
    .ZN(_3115_));
 NOR2_X1 _3860_ (.A1(\fir.p1[4] ),
    .A2(_3115_),
    .ZN(_3116_));
 NAND2_X1 _3861_ (.A1(\fir.p1[4] ),
    .A2(\fir.p1[3] ),
    .ZN(_3117_));
 OR2_X1 _3862_ (.A1(\fir.p1[4] ),
    .A2(\fir.p1[3] ),
    .ZN(_3118_));
 AOI22_X1 _3863_ (.A1(\fir.p1[3] ),
    .A2(\fir.p1[2] ),
    .B1(_3117_),
    .B2(_3118_),
    .ZN(_3119_));
 NOR2_X1 _3864_ (.A1(_3116_),
    .A2(_3119_),
    .ZN(_3120_));
 XNOR2_X1 _3865_ (.A(_3114_),
    .B(_3120_),
    .ZN(_3121_));
 XOR2_X1 _3866_ (.A(_3108_),
    .B(_3121_),
    .Z(_3122_));
 XNOR2_X1 _3867_ (.A(_3107_),
    .B(_3122_),
    .ZN(_3123_));
 XNOR2_X1 _3868_ (.A(_3106_),
    .B(_3123_),
    .ZN(_3124_));
 XNOR2_X1 _3869_ (.A(_3105_),
    .B(_3124_),
    .ZN(_3125_));
 XOR2_X1 _3870_ (.A(_3104_),
    .B(_3125_),
    .Z(_3126_));
 XNOR2_X1 _3871_ (.A(\fir.p2[1] ),
    .B(_3126_),
    .ZN(_3127_));
 XOR2_X1 _3872_ (.A(_3103_),
    .B(_3127_),
    .Z(_3128_));
 XNOR2_X1 _3873_ (.A(\fir.p2[3] ),
    .B(_3128_),
    .ZN(_3129_));
 XNOR2_X1 _3874_ (.A(_3097_),
    .B(_3129_),
    .ZN(_3130_));
 AND2_X1 _3875_ (.A1(_3077_),
    .A2(_3100_),
    .ZN(_3131_));
 INV_X1 _3876_ (.A(_3131_),
    .ZN(_3132_));
 OAI21_X1 _3877_ (.A(_3132_),
    .B1(_3099_),
    .B2(_3078_),
    .ZN(_3133_));
 XOR2_X1 _3878_ (.A(_3130_),
    .B(_3133_),
    .Z(_3134_));
 XNOR2_X1 _3879_ (.A(\fir.p4[4] ),
    .B(_3134_),
    .ZN(_3135_));
 XOR2_X1 _3880_ (.A(_3102_),
    .B(_3135_),
    .Z(_3136_));
 AND2_X1 _3881_ (.A1(\fir.p4[2] ),
    .A2(\fir.p4[1] ),
    .ZN(_3137_));
 OR2_X1 _3882_ (.A1(\fir.p4[0] ),
    .A2(_3137_),
    .ZN(_3138_));
 OAI21_X1 _3883_ (.A(_3138_),
    .B1(\fir.p4[1] ),
    .B2(\fir.p4[2] ),
    .ZN(_3139_));
 OR3_X1 _3884_ (.A1(\fir.p4[2] ),
    .A2(\fir.p4[1] ),
    .A3(\fir.p4[0] ),
    .ZN(_3140_));
 AOI22_X1 _3885_ (.A1(\fir.p4[0] ),
    .A2(_3137_),
    .B1(_3139_),
    .B2(_3140_),
    .ZN(_3141_));
 XNOR2_X1 _3886_ (.A(_3136_),
    .B(_3141_),
    .ZN(_3142_));
 XOR2_X1 _3887_ (.A(\fir.p4[1] ),
    .B(\fir.p4[0] ),
    .Z(_3143_));
 XOR2_X1 _3888_ (.A(_3052_),
    .B(_3076_),
    .Z(_3144_));
 NAND2_X1 _3889_ (.A1(\fir.p4[2] ),
    .A2(_3144_),
    .ZN(_3145_));
 XNOR2_X1 _3890_ (.A(\fir.p4[3] ),
    .B(_3101_),
    .ZN(_3146_));
 XOR2_X1 _3891_ (.A(_3145_),
    .B(_3146_),
    .Z(_3147_));
 AND2_X1 _3892_ (.A1(_3143_),
    .A2(_3147_),
    .ZN(_3148_));
 NOR2_X1 _3893_ (.A1(_3145_),
    .A2(_3146_),
    .ZN(_3149_));
 OAI21_X1 _3894_ (.A(_3142_),
    .B1(_3148_),
    .B2(_3149_),
    .ZN(_3150_));
 NOR2_X1 _3895_ (.A1(_3149_),
    .A2(_3148_),
    .ZN(_3151_));
 XNOR2_X1 _3896_ (.A(_3151_),
    .B(_3142_),
    .ZN(_3152_));
 NAND3_X1 _3897_ (.A1(\fir.p4[1] ),
    .A2(\fir.p4[0] ),
    .A3(_3152_),
    .ZN(_3153_));
 NAND2_X1 _3898_ (.A1(_3150_),
    .A2(_3153_),
    .ZN(_3154_));
 NOR2_X1 _3899_ (.A1(_3102_),
    .A2(_3135_),
    .ZN(_3155_));
 INV_X1 _3900_ (.A(_3141_),
    .ZN(_3156_));
 AOI21_X1 _3901_ (.A(_3155_),
    .B1(_3136_),
    .B2(_3156_),
    .ZN(_3157_));
 NAND2_X1 _3902_ (.A1(\fir.p4[4] ),
    .A2(_3134_),
    .ZN(_3158_));
 NAND2_X1 _3903_ (.A1(_3131_),
    .A2(_3130_),
    .ZN(_3159_));
 NOR2_X1 _3904_ (.A1(_3103_),
    .A2(_3127_),
    .ZN(_3160_));
 AOI21_X1 _3905_ (.A(_3160_),
    .B1(_3128_),
    .B2(\fir.p2[3] ),
    .ZN(_3161_));
 NAND2_X1 _3906_ (.A1(\fir.p2[1] ),
    .A2(_3126_),
    .ZN(_3162_));
 NOR2_X1 _3907_ (.A1(_3104_),
    .A2(_3125_),
    .ZN(_3163_));
 NOR2_X1 _3908_ (.A1(_3105_),
    .A2(_3124_),
    .ZN(_3164_));
 NAND2_X1 _3909_ (.A1(_3106_),
    .A2(_3123_),
    .ZN(_3165_));
 AOI21_X1 _3910_ (.A(_3121_),
    .B1(_3108_),
    .B2(_3107_),
    .ZN(_3166_));
 AOI22_X1 _3911_ (.A1(\fir.p0[4] ),
    .A2(_3109_),
    .B1(_3114_),
    .B2(_3120_),
    .ZN(_3167_));
 AND3_X1 _3912_ (.A1(\fir.p0[3] ),
    .A2(\fir.p0[1] ),
    .A3(_3111_),
    .ZN(_3168_));
 AOI21_X1 _3913_ (.A(_3168_),
    .B1(_3112_),
    .B2(\fir.p0[0] ),
    .ZN(_3169_));
 NAND2_X1 _3914_ (.A1(\fir.p0[4] ),
    .A2(\fir.p0[2] ),
    .ZN(_3170_));
 XOR2_X1 _3915_ (.A(\fir.p0[5] ),
    .B(\fir.p0[3] ),
    .Z(_3171_));
 XNOR2_X1 _3916_ (.A(_3170_),
    .B(_3171_),
    .ZN(_3172_));
 XNOR2_X1 _3917_ (.A(\fir.p0[1] ),
    .B(_3172_),
    .ZN(_3173_));
 XOR2_X1 _3918_ (.A(_3169_),
    .B(_3173_),
    .Z(_3174_));
 NOR2_X1 _3919_ (.A1(\fir.p1[5] ),
    .A2(_3117_),
    .ZN(_3175_));
 OR2_X1 _3920_ (.A1(\fir.p1[5] ),
    .A2(\fir.p1[4] ),
    .ZN(_3176_));
 NAND2_X1 _3921_ (.A1(\fir.p1[5] ),
    .A2(\fir.p1[4] ),
    .ZN(_3177_));
 AOI22_X1 _3922_ (.A1(\fir.p1[4] ),
    .A2(\fir.p1[3] ),
    .B1(_3176_),
    .B2(_3177_),
    .ZN(_3178_));
 NOR2_X1 _3923_ (.A1(_3175_),
    .A2(_3178_),
    .ZN(_3179_));
 XNOR2_X1 _3924_ (.A(_3174_),
    .B(_3179_),
    .ZN(_3180_));
 XNOR2_X1 _3925_ (.A(_3167_),
    .B(_3180_),
    .ZN(_3181_));
 XNOR2_X1 _3926_ (.A(_3116_),
    .B(_3181_),
    .ZN(_3182_));
 XNOR2_X1 _3927_ (.A(_3166_),
    .B(_3182_),
    .ZN(_3183_));
 XOR2_X1 _3928_ (.A(_3165_),
    .B(_3183_),
    .Z(_3184_));
 XNOR2_X1 _3929_ (.A(_3164_),
    .B(_3184_),
    .ZN(_3185_));
 XNOR2_X1 _3930_ (.A(_3163_),
    .B(_3185_),
    .ZN(_3186_));
 XNOR2_X1 _3931_ (.A(\fir.p2[2] ),
    .B(_3186_),
    .ZN(_3187_));
 XOR2_X1 _3932_ (.A(_3162_),
    .B(_3187_),
    .Z(_3188_));
 XOR2_X1 _3933_ (.A(\fir.p2[4] ),
    .B(\fir.p2[0] ),
    .Z(_3189_));
 XNOR2_X1 _3934_ (.A(_3188_),
    .B(_3189_),
    .ZN(_3190_));
 XOR2_X1 _3935_ (.A(_3161_),
    .B(_3190_),
    .Z(_3191_));
 NOR2_X1 _3936_ (.A1(_3096_),
    .A2(_3129_),
    .ZN(_3192_));
 NOR4_X1 _3937_ (.A1(_3078_),
    .A2(_3097_),
    .A3(_3098_),
    .A4(_3129_),
    .ZN(_3193_));
 NOR2_X1 _3938_ (.A1(_3192_),
    .A2(_3193_),
    .ZN(_3194_));
 XNOR2_X1 _3939_ (.A(_3191_),
    .B(_3194_),
    .ZN(_3195_));
 XNOR2_X1 _3940_ (.A(_3159_),
    .B(_3195_),
    .ZN(_3196_));
 XNOR2_X1 _3941_ (.A(\fir.p4[5] ),
    .B(_3196_),
    .ZN(_3197_));
 XOR2_X1 _3942_ (.A(_3158_),
    .B(_3197_),
    .Z(_3198_));
 XOR2_X1 _3943_ (.A(\fir.p4[3] ),
    .B(\fir.p4[2] ),
    .Z(_3199_));
 XNOR2_X1 _3944_ (.A(\fir.p4[1] ),
    .B(_3199_),
    .ZN(_3200_));
 XOR2_X1 _3945_ (.A(_3198_),
    .B(_3200_),
    .Z(_3201_));
 XOR2_X1 _3946_ (.A(_3157_),
    .B(_3201_),
    .Z(_3202_));
 OAI21_X1 _3947_ (.A(\fir.p4[0] ),
    .B1(\fir.p4[1] ),
    .B2(\fir.p4[2] ),
    .ZN(_3203_));
 NAND2_X1 _3948_ (.A1(_3138_),
    .A2(_3203_),
    .ZN(_3204_));
 XOR2_X1 _3949_ (.A(_3202_),
    .B(_3204_),
    .Z(_3205_));
 XNOR2_X1 _3950_ (.A(_3154_),
    .B(_3205_),
    .ZN(_3206_));
 XNOR2_X1 _3951_ (.A(\fir.p3[2] ),
    .B(\fir.p3[0] ),
    .ZN(_3207_));
 XOR2_X1 _3952_ (.A(\fir.p3[1] ),
    .B(_3207_),
    .Z(_3208_));
 INV_X1 _3953_ (.A(_3208_),
    .ZN(_3209_));
 NAND2_X1 _3954_ (.A1(\fir.p3[4] ),
    .A2(_3209_),
    .ZN(_3210_));
 XOR2_X1 _3955_ (.A(\fir.p3[3] ),
    .B(\fir.p3[2] ),
    .Z(_3211_));
 XNOR2_X1 _3956_ (.A(\fir.p3[1] ),
    .B(_3211_),
    .ZN(_3212_));
 XOR2_X1 _3957_ (.A(\fir.p3[5] ),
    .B(_3212_),
    .Z(_3213_));
 XOR2_X1 _3958_ (.A(_3210_),
    .B(_3213_),
    .Z(_3214_));
 XNOR2_X1 _3959_ (.A(_3206_),
    .B(_3214_),
    .ZN(_3215_));
 XOR2_X1 _3960_ (.A(\fir.p3[1] ),
    .B(\fir.p3[0] ),
    .Z(_3216_));
 NAND2_X1 _3961_ (.A1(\fir.p3[3] ),
    .A2(_3216_),
    .ZN(_3217_));
 XNOR2_X1 _3962_ (.A(\fir.p3[4] ),
    .B(_3208_),
    .ZN(_3218_));
 XOR2_X1 _3963_ (.A(_3217_),
    .B(_3218_),
    .Z(_3219_));
 XNOR2_X1 _3964_ (.A(_3143_),
    .B(_3147_),
    .ZN(_3220_));
 INV_X1 _3965_ (.A(net279),
    .ZN(_3221_));
 XNOR2_X1 _3966_ (.A(\fir.p4[2] ),
    .B(_3144_),
    .ZN(_3222_));
 XNOR2_X1 _3967_ (.A(\fir.p2[0] ),
    .B(_3041_),
    .ZN(_3223_));
 OR3_X1 _3968_ (.A1(_3221_),
    .A2(_3222_),
    .A3(_3223_),
    .ZN(_3224_));
 OAI21_X1 _3969_ (.A(_3222_),
    .B1(_3223_),
    .B2(_3221_),
    .ZN(_3225_));
 AND2_X1 _3970_ (.A1(_3224_),
    .A2(_3225_),
    .ZN(_3226_));
 NAND2_X1 _3971_ (.A1(\fir.p4[0] ),
    .A2(_3226_),
    .ZN(_3227_));
 AOI21_X1 _3972_ (.A(_3220_),
    .B1(_3227_),
    .B2(_3224_),
    .ZN(_3228_));
 NAND2_X1 _3973_ (.A1(\fir.p4[1] ),
    .A2(\fir.p4[0] ),
    .ZN(_3229_));
 XNOR2_X1 _3974_ (.A(_3229_),
    .B(_3152_),
    .ZN(_3230_));
 XNOR2_X1 _3975_ (.A(_3228_),
    .B(_3230_),
    .ZN(_3231_));
 OR2_X1 _3976_ (.A1(_3219_),
    .A2(_3231_),
    .ZN(_3232_));
 NAND2_X1 _3977_ (.A1(_3228_),
    .A2(_3230_),
    .ZN(_3233_));
 AOI21_X1 _3978_ (.A(_3215_),
    .B1(_3232_),
    .B2(_3233_),
    .ZN(_3234_));
 XNOR2_X1 _3979_ (.A(\fir.p3[1] ),
    .B(\fir.p3[0] ),
    .ZN(_3235_));
 NAND3_X1 _3980_ (.A1(\fir.p3[3] ),
    .A2(_3216_),
    .A3(_3218_),
    .ZN(_3236_));
 OR3_X1 _3981_ (.A1(_3235_),
    .A2(_3207_),
    .A3(_3236_),
    .ZN(_3237_));
 OAI21_X1 _3982_ (.A(_3236_),
    .B1(_3207_),
    .B2(_3235_),
    .ZN(_3238_));
 NAND2_X1 _3983_ (.A1(_3237_),
    .A2(_3238_),
    .ZN(_3239_));
 NAND2_X1 _3984_ (.A1(_3233_),
    .A2(_3232_),
    .ZN(_3240_));
 XOR2_X1 _3985_ (.A(_3240_),
    .B(_3215_),
    .Z(_3241_));
 NOR2_X1 _3986_ (.A1(_3239_),
    .A2(_3241_),
    .ZN(_3242_));
 NOR2_X1 _3987_ (.A1(_3234_),
    .A2(_3242_),
    .ZN(_3243_));
 AOI21_X1 _3988_ (.A(_3205_),
    .B1(_3153_),
    .B2(_3150_),
    .ZN(_3244_));
 AOI21_X1 _3989_ (.A(_3244_),
    .B1(_3206_),
    .B2(_3214_),
    .ZN(_3245_));
 NAND3_X1 _3990_ (.A1(_3138_),
    .A2(_3202_),
    .A3(_3203_),
    .ZN(_3246_));
 OAI21_X1 _3991_ (.A(_3246_),
    .B1(_3201_),
    .B2(_3157_),
    .ZN(_3247_));
 NOR2_X1 _3992_ (.A1(_3158_),
    .A2(_3197_),
    .ZN(_3248_));
 INV_X1 _3993_ (.A(_3198_),
    .ZN(_3249_));
 NOR2_X1 _3994_ (.A1(_3249_),
    .A2(_3200_),
    .ZN(_3250_));
 NOR2_X1 _3995_ (.A1(_3248_),
    .A2(_3250_),
    .ZN(_3251_));
 NAND2_X1 _3996_ (.A1(\fir.p4[5] ),
    .A2(_3196_),
    .ZN(_3252_));
 NAND2_X1 _3997_ (.A1(_3193_),
    .A2(_3191_),
    .ZN(_3253_));
 NAND3_X1 _3998_ (.A1(_3131_),
    .A2(_3130_),
    .A3(_3195_),
    .ZN(_3254_));
 NAND2_X1 _3999_ (.A1(_3253_),
    .A2(_3254_),
    .ZN(_3255_));
 NAND2_X1 _4000_ (.A1(\fir.p2[4] ),
    .A2(\fir.p2[0] ),
    .ZN(_3256_));
 NOR2_X1 _4001_ (.A1(_3162_),
    .A2(_3187_),
    .ZN(_3257_));
 AOI21_X1 _4002_ (.A(_3257_),
    .B1(_3188_),
    .B2(_3189_),
    .ZN(_3258_));
 NAND2_X1 _4003_ (.A1(\fir.p2[2] ),
    .A2(_3186_),
    .ZN(_3259_));
 NOR2_X1 _4004_ (.A1(_3165_),
    .A2(_3183_),
    .ZN(_3260_));
 NAND2_X1 _4005_ (.A1(_3166_),
    .A2(_3182_),
    .ZN(_3261_));
 NOR2_X1 _4006_ (.A1(_3167_),
    .A2(_3180_),
    .ZN(_3262_));
 NAND2_X1 _4007_ (.A1(_3167_),
    .A2(_3180_),
    .ZN(_3263_));
 AOI21_X1 _4008_ (.A(_3262_),
    .B1(_3263_),
    .B2(_3116_),
    .ZN(_3264_));
 NOR2_X1 _4009_ (.A1(_3169_),
    .A2(_3173_),
    .ZN(_3265_));
 AOI21_X1 _4010_ (.A(_3265_),
    .B1(_3174_),
    .B2(_3179_),
    .ZN(_3266_));
 AND3_X1 _4011_ (.A1(\fir.p0[4] ),
    .A2(\fir.p0[2] ),
    .A3(_3171_),
    .ZN(_3267_));
 AOI21_X1 _4012_ (.A(_3267_),
    .B1(_3172_),
    .B2(\fir.p0[1] ),
    .ZN(_3268_));
 NAND2_X1 _4013_ (.A1(\fir.p0[5] ),
    .A2(\fir.p0[3] ),
    .ZN(_3269_));
 XOR2_X1 _4014_ (.A(\fir.p0[6] ),
    .B(\fir.p0[4] ),
    .Z(_3270_));
 XNOR2_X1 _4015_ (.A(_3269_),
    .B(_3270_),
    .ZN(_3271_));
 XNOR2_X1 _4016_ (.A(\fir.p0[2] ),
    .B(_3271_),
    .ZN(_3272_));
 XOR2_X1 _4017_ (.A(_3268_),
    .B(_3272_),
    .Z(_3273_));
 NOR2_X1 _4018_ (.A1(\fir.p1[6] ),
    .A2(_3177_),
    .ZN(_3274_));
 OR2_X1 _4019_ (.A1(\fir.p1[6] ),
    .A2(\fir.p1[5] ),
    .ZN(_3275_));
 NAND2_X1 _4020_ (.A1(\fir.p1[6] ),
    .A2(\fir.p1[5] ),
    .ZN(_3276_));
 AOI22_X1 _4021_ (.A1(\fir.p1[5] ),
    .A2(\fir.p1[4] ),
    .B1(_3275_),
    .B2(_3276_),
    .ZN(_3277_));
 NOR2_X1 _4022_ (.A1(_3274_),
    .A2(_3277_),
    .ZN(_3278_));
 XOR2_X1 _4023_ (.A(_3273_),
    .B(_3278_),
    .Z(_3279_));
 XNOR2_X1 _4024_ (.A(_3266_),
    .B(_3279_),
    .ZN(_3280_));
 XNOR2_X1 _4025_ (.A(_0004_),
    .B(_3175_),
    .ZN(_3281_));
 XNOR2_X1 _4026_ (.A(_3280_),
    .B(_3281_),
    .ZN(_3282_));
 XOR2_X1 _4027_ (.A(_3264_),
    .B(_3282_),
    .Z(_3283_));
 XNOR2_X1 _4028_ (.A(_3261_),
    .B(_3283_),
    .ZN(_3284_));
 XOR2_X1 _4029_ (.A(_3260_),
    .B(_3284_),
    .Z(_3285_));
 AND2_X1 _4030_ (.A1(_3105_),
    .A2(_3124_),
    .ZN(_3286_));
 XNOR2_X1 _4031_ (.A(_3165_),
    .B(_3183_),
    .ZN(_3287_));
 NOR4_X1 _4032_ (.A1(_3104_),
    .A2(_3164_),
    .A3(_3286_),
    .A4(_3287_),
    .ZN(_3288_));
 AND2_X1 _4033_ (.A1(_3164_),
    .A2(_3184_),
    .ZN(_3289_));
 OAI21_X1 _4034_ (.A(_3285_),
    .B1(_3288_),
    .B2(_3289_),
    .ZN(_3290_));
 OR3_X1 _4035_ (.A1(_3289_),
    .A2(_3288_),
    .A3(_3285_),
    .ZN(_3291_));
 AND2_X1 _4036_ (.A1(_3290_),
    .A2(_3291_),
    .ZN(_3292_));
 XNOR2_X1 _4037_ (.A(\fir.p2[3] ),
    .B(_3292_),
    .ZN(_3293_));
 XOR2_X1 _4038_ (.A(_3259_),
    .B(_3293_),
    .Z(_3294_));
 XOR2_X1 _4039_ (.A(\fir.p2[5] ),
    .B(\fir.p2[1] ),
    .Z(_3295_));
 XNOR2_X1 _4040_ (.A(_3294_),
    .B(_3295_),
    .ZN(_3296_));
 XOR2_X1 _4041_ (.A(_3258_),
    .B(_3296_),
    .Z(_3297_));
 XNOR2_X1 _4042_ (.A(_3256_),
    .B(_3297_),
    .ZN(_3298_));
 NOR2_X1 _4043_ (.A1(_3161_),
    .A2(_3190_),
    .ZN(_3299_));
 AND2_X1 _4044_ (.A1(_3192_),
    .A2(_3191_),
    .ZN(_3300_));
 NOR2_X1 _4045_ (.A1(_3299_),
    .A2(_3300_),
    .ZN(_3301_));
 XNOR2_X1 _4046_ (.A(_3298_),
    .B(_3301_),
    .ZN(_3302_));
 XOR2_X1 _4047_ (.A(_3255_),
    .B(_3302_),
    .Z(_3303_));
 XNOR2_X1 _4048_ (.A(\fir.p4[6] ),
    .B(_3303_),
    .ZN(_3304_));
 XOR2_X1 _4049_ (.A(_3252_),
    .B(_3304_),
    .Z(_3305_));
 XOR2_X1 _4050_ (.A(\fir.p4[4] ),
    .B(\fir.p4[3] ),
    .Z(_3306_));
 XNOR2_X1 _4051_ (.A(\fir.p4[2] ),
    .B(_3306_),
    .ZN(_3307_));
 XNOR2_X1 _4052_ (.A(_3305_),
    .B(_3307_),
    .ZN(_3308_));
 XNOR2_X1 _4053_ (.A(_3251_),
    .B(_3308_),
    .ZN(_3309_));
 AND2_X1 _4054_ (.A1(\fir.p4[3] ),
    .A2(\fir.p4[2] ),
    .ZN(_3310_));
 AOI21_X1 _4055_ (.A(_3310_),
    .B1(_3199_),
    .B2(\fir.p4[1] ),
    .ZN(_3311_));
 XNOR2_X1 _4056_ (.A(_3143_),
    .B(_3311_),
    .ZN(_3312_));
 XOR2_X1 _4057_ (.A(_3309_),
    .B(_3312_),
    .Z(_3313_));
 XNOR2_X1 _4058_ (.A(_3247_),
    .B(_3313_),
    .ZN(_3314_));
 INV_X1 _4059_ (.A(_3212_),
    .ZN(_3315_));
 NAND2_X1 _4060_ (.A1(\fir.p3[5] ),
    .A2(_3315_),
    .ZN(_3316_));
 XOR2_X1 _4061_ (.A(\fir.p3[4] ),
    .B(\fir.p3[3] ),
    .Z(_3317_));
 XNOR2_X1 _4062_ (.A(\fir.p3[2] ),
    .B(_3317_),
    .ZN(_3318_));
 XOR2_X1 _4063_ (.A(\fir.p3[6] ),
    .B(_3318_),
    .Z(_3319_));
 XOR2_X1 _4064_ (.A(_3203_),
    .B(_3319_),
    .Z(_3320_));
 XNOR2_X1 _4065_ (.A(_3316_),
    .B(_3320_),
    .ZN(_3321_));
 INV_X1 _4066_ (.A(_3321_),
    .ZN(_3322_));
 XNOR2_X1 _4067_ (.A(_3314_),
    .B(_3322_),
    .ZN(_3323_));
 XOR2_X1 _4068_ (.A(_3245_),
    .B(_3323_),
    .Z(_3324_));
 NOR2_X1 _4069_ (.A1(_3210_),
    .A2(_3213_),
    .ZN(_3325_));
 AOI21_X1 _4070_ (.A(\fir.p3[1] ),
    .B1(\fir.p3[0] ),
    .B2(\fir.p3[2] ),
    .ZN(_3326_));
 INV_X1 _4071_ (.A(_3326_),
    .ZN(_3327_));
 NAND2_X1 _4072_ (.A1(\fir.p3[0] ),
    .A2(_3327_),
    .ZN(_3328_));
 AND2_X1 _4073_ (.A1(\fir.p3[3] ),
    .A2(\fir.p3[2] ),
    .ZN(_3329_));
 AOI21_X1 _4074_ (.A(_3329_),
    .B1(_3211_),
    .B2(\fir.p3[1] ),
    .ZN(_3330_));
 XNOR2_X1 _4075_ (.A(_3216_),
    .B(_3330_),
    .ZN(_3331_));
 XNOR2_X1 _4076_ (.A(_3328_),
    .B(_3331_),
    .ZN(_3332_));
 XOR2_X1 _4077_ (.A(_3325_),
    .B(_3332_),
    .Z(_3333_));
 XNOR2_X1 _4078_ (.A(_3324_),
    .B(_3333_),
    .ZN(_3334_));
 NOR2_X1 _4079_ (.A1(_3243_),
    .A2(_3334_),
    .ZN(_3335_));
 XNOR2_X1 _4080_ (.A(_3243_),
    .B(_3334_),
    .ZN(_3336_));
 NOR2_X1 _4081_ (.A1(_3237_),
    .A2(_3336_),
    .ZN(_3337_));
 NOR2_X1 _4082_ (.A1(_3335_),
    .A2(_3337_),
    .ZN(_3338_));
 AND2_X1 _4083_ (.A1(_3325_),
    .A2(_3332_),
    .ZN(_3339_));
 OR2_X1 _4084_ (.A1(_3245_),
    .A2(_3323_),
    .ZN(_3340_));
 NAND2_X1 _4085_ (.A1(_3324_),
    .A2(_3333_),
    .ZN(_3341_));
 NAND2_X1 _4086_ (.A1(_3340_),
    .A2(_3341_),
    .ZN(_3342_));
 NOR2_X1 _4087_ (.A1(_3314_),
    .A2(_3322_),
    .ZN(_3343_));
 AOI21_X1 _4088_ (.A(_3343_),
    .B1(_3313_),
    .B2(_3247_),
    .ZN(_3344_));
 OAI21_X1 _4089_ (.A(_3308_),
    .B1(_3250_),
    .B2(_3248_),
    .ZN(_3345_));
 NAND2_X1 _4090_ (.A1(_3309_),
    .A2(_3312_),
    .ZN(_3346_));
 NAND2_X1 _4091_ (.A1(_3345_),
    .A2(_3346_),
    .ZN(_3347_));
 NOR2_X1 _4092_ (.A1(_3252_),
    .A2(_3304_),
    .ZN(_3348_));
 INV_X1 _4093_ (.A(_3307_),
    .ZN(_3349_));
 AOI21_X1 _4094_ (.A(_3348_),
    .B1(_3305_),
    .B2(_3349_),
    .ZN(_3350_));
 NAND2_X1 _4095_ (.A1(\fir.p4[6] ),
    .A2(_3303_),
    .ZN(_3351_));
 AOI22_X1 _4096_ (.A1(_3300_),
    .A2(_3298_),
    .B1(_3302_),
    .B2(_3255_),
    .ZN(_3352_));
 NAND2_X1 _4097_ (.A1(_3299_),
    .A2(_3298_),
    .ZN(_3353_));
 NAND3_X1 _4098_ (.A1(\fir.p2[4] ),
    .A2(\fir.p2[0] ),
    .A3(_3297_),
    .ZN(_3354_));
 OAI21_X1 _4099_ (.A(_3354_),
    .B1(_3296_),
    .B2(_3258_),
    .ZN(_3355_));
 NOR2_X1 _4100_ (.A1(_3259_),
    .A2(_3293_),
    .ZN(_3356_));
 AOI21_X1 _4101_ (.A(_3356_),
    .B1(_3294_),
    .B2(_3295_),
    .ZN(_3357_));
 NAND2_X1 _4102_ (.A1(\fir.p2[3] ),
    .A2(_3292_),
    .ZN(_3358_));
 AND3_X1 _4103_ (.A1(_3166_),
    .A2(_3182_),
    .A3(_3283_),
    .ZN(_3359_));
 NOR2_X1 _4104_ (.A1(_3264_),
    .A2(_3282_),
    .ZN(_3360_));
 NOR3_X1 _4105_ (.A1(\fir.p1[5] ),
    .A2(_0004_),
    .A3(_3117_),
    .ZN(_3361_));
 NAND2_X1 _4106_ (.A1(_3174_),
    .A2(_3179_),
    .ZN(_3362_));
 OAI21_X1 _4107_ (.A(_3362_),
    .B1(_3173_),
    .B2(_3169_),
    .ZN(_3363_));
 AOI22_X1 _4108_ (.A1(_3363_),
    .A2(_3279_),
    .B1(_3280_),
    .B2(_3281_),
    .ZN(_3364_));
 NOR2_X1 _4109_ (.A1(_3268_),
    .A2(_3272_),
    .ZN(_3365_));
 AOI21_X1 _4110_ (.A(_3365_),
    .B1(_3273_),
    .B2(_3278_),
    .ZN(_3366_));
 AND3_X1 _4111_ (.A1(\fir.p0[5] ),
    .A2(\fir.p0[3] ),
    .A3(_3270_),
    .ZN(_3367_));
 AOI21_X1 _4112_ (.A(_3367_),
    .B1(_3271_),
    .B2(\fir.p0[2] ),
    .ZN(_3368_));
 NAND2_X1 _4113_ (.A1(\fir.p0[6] ),
    .A2(\fir.p0[4] ),
    .ZN(_3369_));
 XOR2_X1 _4114_ (.A(\fir.p0[7] ),
    .B(\fir.p0[5] ),
    .Z(_3370_));
 XNOR2_X1 _4115_ (.A(_3369_),
    .B(_3370_),
    .ZN(_3371_));
 XNOR2_X1 _4116_ (.A(\fir.p0[3] ),
    .B(_3371_),
    .ZN(_3372_));
 XOR2_X1 _4117_ (.A(_3368_),
    .B(_3372_),
    .Z(_3373_));
 OR2_X1 _4118_ (.A1(\fir.p1[7] ),
    .A2(\fir.p1[6] ),
    .ZN(_3374_));
 NAND2_X1 _4119_ (.A1(\fir.p1[7] ),
    .A2(\fir.p1[6] ),
    .ZN(_3375_));
 AOI22_X1 _4120_ (.A1(\fir.p1[6] ),
    .A2(\fir.p1[5] ),
    .B1(_3374_),
    .B2(_3375_),
    .ZN(_3376_));
 NOR2_X1 _4121_ (.A1(\fir.p1[7] ),
    .A2(_3276_),
    .ZN(_3377_));
 NOR2_X1 _4122_ (.A1(_3376_),
    .A2(_3377_),
    .ZN(_3378_));
 XNOR2_X1 _4123_ (.A(_3373_),
    .B(_3378_),
    .ZN(_3379_));
 XOR2_X1 _4124_ (.A(_3366_),
    .B(_3379_),
    .Z(_3380_));
 XNOR2_X1 _4125_ (.A(_0003_),
    .B(_3274_),
    .ZN(_3381_));
 XNOR2_X1 _4126_ (.A(_3380_),
    .B(_3381_),
    .ZN(_3382_));
 XOR2_X1 _4127_ (.A(_3364_),
    .B(_3382_),
    .Z(_3383_));
 XOR2_X1 _4128_ (.A(_3361_),
    .B(_3383_),
    .Z(_3384_));
 XOR2_X1 _4129_ (.A(_3360_),
    .B(_3384_),
    .Z(_3385_));
 XNOR2_X1 _4130_ (.A(_3359_),
    .B(_3385_),
    .ZN(_3386_));
 NAND2_X1 _4131_ (.A1(_3260_),
    .A2(_3284_),
    .ZN(_3387_));
 NAND2_X1 _4132_ (.A1(_3387_),
    .A2(_3290_),
    .ZN(_3388_));
 XNOR2_X1 _4133_ (.A(_3386_),
    .B(_3388_),
    .ZN(_3389_));
 XNOR2_X1 _4134_ (.A(\fir.p2[4] ),
    .B(_3389_),
    .ZN(_3390_));
 XOR2_X1 _4135_ (.A(_3358_),
    .B(_3390_),
    .Z(_3391_));
 XOR2_X1 _4136_ (.A(\fir.p2[6] ),
    .B(\fir.p2[2] ),
    .Z(_3392_));
 XNOR2_X1 _4137_ (.A(_3391_),
    .B(_3392_),
    .ZN(_3393_));
 XOR2_X1 _4138_ (.A(_3357_),
    .B(_3393_),
    .Z(_3394_));
 NAND2_X1 _4139_ (.A1(\fir.p2[5] ),
    .A2(\fir.p2[1] ),
    .ZN(_3395_));
 XOR2_X1 _4140_ (.A(_0009_),
    .B(_3395_),
    .Z(_3396_));
 XNOR2_X1 _4141_ (.A(_3394_),
    .B(_3396_),
    .ZN(_3397_));
 XOR2_X1 _4142_ (.A(_3355_),
    .B(_3397_),
    .Z(_3398_));
 XNOR2_X1 _4143_ (.A(_3353_),
    .B(_3398_),
    .ZN(_3399_));
 XOR2_X1 _4144_ (.A(_3352_),
    .B(_3399_),
    .Z(_3400_));
 XNOR2_X1 _4145_ (.A(\fir.p4[7] ),
    .B(_3400_),
    .ZN(_3401_));
 XOR2_X1 _4146_ (.A(_3351_),
    .B(_3401_),
    .Z(_3402_));
 XOR2_X1 _4147_ (.A(\fir.p4[5] ),
    .B(\fir.p4[4] ),
    .Z(_3403_));
 XNOR2_X1 _4148_ (.A(\fir.p4[3] ),
    .B(_3403_),
    .ZN(_3404_));
 INV_X1 _4149_ (.A(_3404_),
    .ZN(_3405_));
 XNOR2_X1 _4150_ (.A(_3402_),
    .B(_3405_),
    .ZN(_3406_));
 XOR2_X1 _4151_ (.A(_3350_),
    .B(_3406_),
    .Z(_3407_));
 AND2_X1 _4152_ (.A1(\fir.p4[4] ),
    .A2(\fir.p4[3] ),
    .ZN(_3408_));
 AOI21_X1 _4153_ (.A(_3408_),
    .B1(_3306_),
    .B2(\fir.p4[2] ),
    .ZN(_3409_));
 XNOR2_X1 _4154_ (.A(_3141_),
    .B(_3409_),
    .ZN(_3410_));
 XOR2_X1 _4155_ (.A(_3229_),
    .B(_3410_),
    .Z(_3411_));
 XNOR2_X1 _4156_ (.A(_3407_),
    .B(_3411_),
    .ZN(_3412_));
 XNOR2_X1 _4157_ (.A(_3347_),
    .B(_3412_),
    .ZN(_3413_));
 INV_X1 _4158_ (.A(_3318_),
    .ZN(_3414_));
 NAND2_X1 _4159_ (.A1(\fir.p3[6] ),
    .A2(_3414_),
    .ZN(_3415_));
 XNOR2_X1 _4160_ (.A(\fir.p4[1] ),
    .B(\fir.p4[0] ),
    .ZN(_3416_));
 NOR2_X1 _4161_ (.A1(_3416_),
    .A2(_3311_),
    .ZN(_3417_));
 XOR2_X1 _4162_ (.A(\fir.p3[5] ),
    .B(\fir.p3[4] ),
    .Z(_3418_));
 XNOR2_X1 _4163_ (.A(\fir.p3[3] ),
    .B(_3418_),
    .ZN(_3419_));
 XOR2_X1 _4164_ (.A(\fir.p3[7] ),
    .B(_3419_),
    .Z(_3420_));
 XOR2_X1 _4165_ (.A(_3417_),
    .B(_3420_),
    .Z(_3421_));
 XOR2_X1 _4166_ (.A(_3415_),
    .B(_3421_),
    .Z(_3422_));
 XNOR2_X1 _4167_ (.A(_3413_),
    .B(_3422_),
    .ZN(_3423_));
 XOR2_X1 _4168_ (.A(_3344_),
    .B(_3423_),
    .Z(_3424_));
 NAND3_X1 _4169_ (.A1(\fir.p3[0] ),
    .A2(_3327_),
    .A3(_3331_),
    .ZN(_3425_));
 NOR2_X1 _4170_ (.A1(_3235_),
    .A2(_3330_),
    .ZN(_3426_));
 NAND2_X1 _4171_ (.A1(\fir.p3[1] ),
    .A2(\fir.p3[0] ),
    .ZN(_3427_));
 AND2_X1 _4172_ (.A1(\fir.p3[4] ),
    .A2(\fir.p3[3] ),
    .ZN(_3428_));
 AOI21_X1 _4173_ (.A(_3428_),
    .B1(_3317_),
    .B2(\fir.p3[2] ),
    .ZN(_3429_));
 XNOR2_X1 _4174_ (.A(_3208_),
    .B(_3429_),
    .ZN(_3430_));
 XOR2_X1 _4175_ (.A(_3427_),
    .B(_3430_),
    .Z(_3431_));
 XNOR2_X1 _4176_ (.A(_3426_),
    .B(_3431_),
    .ZN(_3432_));
 NAND3_X1 _4177_ (.A1(\fir.p3[5] ),
    .A2(_3315_),
    .A3(_3320_),
    .ZN(_3433_));
 OR2_X1 _4178_ (.A1(_3203_),
    .A2(_3319_),
    .ZN(_3434_));
 AOI21_X1 _4179_ (.A(_3432_),
    .B1(_3433_),
    .B2(_3434_),
    .ZN(_3435_));
 INV_X1 _4180_ (.A(_3435_),
    .ZN(_3436_));
 NAND3_X1 _4181_ (.A1(_3434_),
    .A2(_3433_),
    .A3(_3432_),
    .ZN(_3437_));
 NAND2_X1 _4182_ (.A1(_3436_),
    .A2(_3437_),
    .ZN(_3438_));
 XOR2_X1 _4183_ (.A(_3425_),
    .B(_3438_),
    .Z(_3439_));
 XNOR2_X1 _4184_ (.A(_3424_),
    .B(_3439_),
    .ZN(_3440_));
 XNOR2_X1 _4185_ (.A(_3342_),
    .B(_3440_),
    .ZN(_3441_));
 XNOR2_X1 _4186_ (.A(_3339_),
    .B(_3441_),
    .ZN(_3442_));
 NOR2_X1 _4187_ (.A1(_3338_),
    .A2(_3442_),
    .ZN(_3443_));
 XNOR2_X1 _4188_ (.A(_3219_),
    .B(_3231_),
    .ZN(_3444_));
 AND3_X1 _4189_ (.A1(_3224_),
    .A2(_3227_),
    .A3(_3220_),
    .ZN(_3445_));
 NOR2_X1 _4190_ (.A1(_3228_),
    .A2(_3445_),
    .ZN(_3446_));
 XOR2_X1 _4191_ (.A(\fir.p1[0] ),
    .B(\fir.p0[0] ),
    .Z(_3447_));
 NAND2_X1 _4192_ (.A1(\fir.p4[0] ),
    .A2(_3447_),
    .ZN(_3448_));
 XNOR2_X1 _4193_ (.A(_3221_),
    .B(_3223_),
    .ZN(_3449_));
 XNOR2_X1 _4194_ (.A(\fir.p4[0] ),
    .B(_3226_),
    .ZN(_3450_));
 NOR3_X1 _4195_ (.A1(_3448_),
    .A2(_3449_),
    .A3(_3450_),
    .ZN(_3451_));
 XNOR2_X1 _4196_ (.A(_3446_),
    .B(_3451_),
    .ZN(_3452_));
 NAND2_X1 _4197_ (.A1(\fir.p3[2] ),
    .A2(\fir.p3[0] ),
    .ZN(_3453_));
 XNOR2_X1 _4198_ (.A(\fir.p3[3] ),
    .B(_3216_),
    .ZN(_3454_));
 XNOR2_X1 _4199_ (.A(_3453_),
    .B(_3454_),
    .ZN(_3455_));
 OR2_X1 _4200_ (.A1(_3452_),
    .A2(_3455_),
    .ZN(_3456_));
 NAND2_X1 _4201_ (.A1(_3446_),
    .A2(_3451_),
    .ZN(_3457_));
 AOI21_X1 _4202_ (.A(_3444_),
    .B1(_3456_),
    .B2(_3457_),
    .ZN(_3458_));
 NAND2_X1 _4203_ (.A1(_3457_),
    .A2(_3456_),
    .ZN(_3459_));
 XOR2_X1 _4204_ (.A(_3459_),
    .B(_3444_),
    .Z(_3460_));
 NOR3_X1 _4205_ (.A1(_3329_),
    .A2(_3328_),
    .A3(_3460_),
    .ZN(_3461_));
 NOR2_X1 _4206_ (.A1(_3458_),
    .A2(_3461_),
    .ZN(_3462_));
 XNOR2_X1 _4207_ (.A(_3239_),
    .B(_3241_),
    .ZN(_3463_));
 XNOR2_X1 _4208_ (.A(_3462_),
    .B(_3463_),
    .ZN(_3464_));
 NAND3_X1 _4209_ (.A1(\fir.p3[1] ),
    .A2(\fir.p3[0] ),
    .A3(_3329_),
    .ZN(_3465_));
 OAI22_X1 _4210_ (.A1(_3462_),
    .A2(_3463_),
    .B1(_3464_),
    .B2(_3465_),
    .ZN(_3466_));
 XOR2_X1 _4211_ (.A(_3237_),
    .B(_3336_),
    .Z(_3467_));
 AND2_X1 _4212_ (.A1(_3466_),
    .A2(_3467_),
    .ZN(_3468_));
 XNOR2_X1 _4213_ (.A(_3466_),
    .B(_3467_),
    .ZN(_3469_));
 XOR2_X1 _4214_ (.A(_3465_),
    .B(_3464_),
    .Z(_3470_));
 NOR2_X1 _4215_ (.A1(_3448_),
    .A2(_3449_),
    .ZN(_3471_));
 XOR2_X1 _4216_ (.A(_3471_),
    .B(_3450_),
    .Z(_3472_));
 NOR2_X1 _4217_ (.A1(_3207_),
    .A2(_3472_),
    .ZN(_3473_));
 XOR2_X1 _4218_ (.A(_3452_),
    .B(_3455_),
    .Z(_3474_));
 NOR2_X1 _4219_ (.A1(_3329_),
    .A2(_3328_),
    .ZN(_3475_));
 XNOR2_X1 _4220_ (.A(_3475_),
    .B(_3460_),
    .ZN(_3476_));
 NAND3_X1 _4221_ (.A1(_3473_),
    .A2(_3474_),
    .A3(_3476_),
    .ZN(_3477_));
 INV_X1 _4222_ (.A(_3477_),
    .ZN(_3478_));
 NAND2_X1 _4223_ (.A1(_3470_),
    .A2(_3478_),
    .ZN(_3479_));
 XNOR2_X1 _4224_ (.A(_3470_),
    .B(_3478_),
    .ZN(_3480_));
 INV_X1 _4225_ (.A(_3480_),
    .ZN(_3481_));
 AOI21_X1 _4226_ (.A(_3476_),
    .B1(_3474_),
    .B2(_3473_),
    .ZN(_3482_));
 NOR2_X1 _4227_ (.A1(_3478_),
    .A2(_3482_),
    .ZN(_3483_));
 XOR2_X1 _4228_ (.A(_3448_),
    .B(_3449_),
    .Z(_3484_));
 NAND2_X1 _4229_ (.A1(\fir.p3[1] ),
    .A2(_3484_),
    .ZN(_3485_));
 XNOR2_X1 _4230_ (.A(_3207_),
    .B(_3472_),
    .ZN(_3486_));
 NOR2_X1 _4231_ (.A1(_3485_),
    .A2(_3486_),
    .ZN(_3487_));
 XOR2_X1 _4232_ (.A(_3473_),
    .B(_3474_),
    .Z(_3488_));
 NAND3_X1 _4233_ (.A1(_3483_),
    .A2(_3487_),
    .A3(_3488_),
    .ZN(_3489_));
 XNOR2_X1 _4234_ (.A(\fir.p4[0] ),
    .B(_3447_),
    .ZN(_3490_));
 INV_X1 _4235_ (.A(_3490_),
    .ZN(_3491_));
 NAND2_X1 _4236_ (.A1(\fir.p3[0] ),
    .A2(_3491_),
    .ZN(_3492_));
 XNOR2_X1 _4237_ (.A(\fir.p3[1] ),
    .B(_3484_),
    .ZN(_3493_));
 NOR2_X1 _4238_ (.A1(_3492_),
    .A2(_3493_),
    .ZN(_3494_));
 XOR2_X1 _4239_ (.A(_3485_),
    .B(_3486_),
    .Z(_3495_));
 AND2_X1 _4240_ (.A1(_3494_),
    .A2(_3495_),
    .ZN(_3496_));
 NAND2_X1 _4241_ (.A1(_3488_),
    .A2(_3496_),
    .ZN(_3497_));
 NAND2_X1 _4242_ (.A1(_3487_),
    .A2(_3488_),
    .ZN(_3498_));
 XOR2_X1 _4243_ (.A(_3483_),
    .B(_3498_),
    .Z(_3499_));
 OAI21_X1 _4244_ (.A(_3489_),
    .B1(_3497_),
    .B2(_3499_),
    .ZN(_3500_));
 NAND2_X1 _4245_ (.A1(_3481_),
    .A2(_3500_),
    .ZN(_3501_));
 AOI21_X1 _4246_ (.A(_3469_),
    .B1(_3479_),
    .B2(_3501_),
    .ZN(_3502_));
 OR2_X1 _4247_ (.A1(_3468_),
    .A2(_3502_),
    .ZN(_3503_));
 XOR2_X1 _4248_ (.A(_3338_),
    .B(_3442_),
    .Z(_3504_));
 AOI21_X1 _4249_ (.A(_3443_),
    .B1(_3503_),
    .B2(_3504_),
    .ZN(_3505_));
 AOI21_X1 _4250_ (.A(_3440_),
    .B1(_3341_),
    .B2(_3340_),
    .ZN(_3506_));
 AOI21_X1 _4251_ (.A(_3506_),
    .B1(_3441_),
    .B2(_3339_),
    .ZN(_3507_));
 NOR2_X1 _4252_ (.A1(_3344_),
    .A2(_3423_),
    .ZN(_3508_));
 AOI21_X1 _4253_ (.A(_3508_),
    .B1(_3424_),
    .B2(_3439_),
    .ZN(_3509_));
 AOI21_X1 _4254_ (.A(_3412_),
    .B1(_3346_),
    .B2(_3345_),
    .ZN(_3510_));
 AOI21_X1 _4255_ (.A(_3510_),
    .B1(_3413_),
    .B2(_3422_),
    .ZN(_3511_));
 NOR2_X1 _4256_ (.A1(_3350_),
    .A2(_3406_),
    .ZN(_3512_));
 AOI21_X1 _4257_ (.A(_3512_),
    .B1(_3407_),
    .B2(_3411_),
    .ZN(_3513_));
 NOR2_X1 _4258_ (.A1(_3351_),
    .A2(_3401_),
    .ZN(_3514_));
 AOI21_X1 _4259_ (.A(_3514_),
    .B1(_3402_),
    .B2(_3405_),
    .ZN(_3515_));
 NAND2_X1 _4260_ (.A1(\fir.p4[7] ),
    .A2(_3400_),
    .ZN(_3516_));
 INV_X1 _4261_ (.A(net267),
    .ZN(_3517_));
 OAI22_X1 _4262_ (.A1(_3353_),
    .A2(_3398_),
    .B1(_3399_),
    .B2(_3352_),
    .ZN(_3518_));
 INV_X1 _4263_ (.A(_3355_),
    .ZN(_3519_));
 NOR2_X1 _4264_ (.A1(_3519_),
    .A2(_3397_),
    .ZN(_3520_));
 NOR2_X1 _4265_ (.A1(_0009_),
    .A2(_3395_),
    .ZN(_3521_));
 NOR2_X1 _4266_ (.A1(_3357_),
    .A2(_3393_),
    .ZN(_3522_));
 AOI21_X1 _4267_ (.A(_3522_),
    .B1(_3394_),
    .B2(_3396_),
    .ZN(_3523_));
 NOR2_X1 _4268_ (.A1(_3358_),
    .A2(_3390_),
    .ZN(_3524_));
 AOI21_X1 _4269_ (.A(_3524_),
    .B1(_3391_),
    .B2(_3392_),
    .ZN(_3525_));
 NAND2_X1 _4270_ (.A1(\fir.p2[4] ),
    .A2(_3389_),
    .ZN(_3526_));
 AND2_X1 _4271_ (.A1(_3260_),
    .A2(_3284_),
    .ZN(_3527_));
 OAI21_X1 _4272_ (.A(_3385_),
    .B1(_3527_),
    .B2(_3359_),
    .ZN(_3528_));
 OAI21_X1 _4273_ (.A(_3528_),
    .B1(_3386_),
    .B2(_3290_),
    .ZN(_3529_));
 AND2_X1 _4274_ (.A1(_3360_),
    .A2(_3384_),
    .ZN(_3530_));
 NOR2_X1 _4275_ (.A1(_3364_),
    .A2(_3382_),
    .ZN(_3531_));
 AOI21_X1 _4276_ (.A(_3531_),
    .B1(_3383_),
    .B2(_3361_),
    .ZN(_3532_));
 NOR3_X1 _4277_ (.A1(\fir.p1[6] ),
    .A2(_0003_),
    .A3(_3177_),
    .ZN(_3533_));
 NOR2_X1 _4278_ (.A1(_3366_),
    .A2(_3379_),
    .ZN(_3534_));
 AOI21_X1 _4279_ (.A(_3534_),
    .B1(_3380_),
    .B2(_3381_),
    .ZN(_3535_));
 NOR2_X1 _4280_ (.A1(_3368_),
    .A2(_3372_),
    .ZN(_3536_));
 AOI21_X1 _4281_ (.A(_3536_),
    .B1(_3373_),
    .B2(_3378_),
    .ZN(_3537_));
 AND3_X1 _4282_ (.A1(\fir.p0[6] ),
    .A2(\fir.p0[4] ),
    .A3(_3370_),
    .ZN(_3538_));
 AOI21_X1 _4283_ (.A(_3538_),
    .B1(_3371_),
    .B2(\fir.p0[3] ),
    .ZN(_3539_));
 NAND2_X1 _4284_ (.A1(\fir.p0[7] ),
    .A2(\fir.p0[5] ),
    .ZN(_3540_));
 XOR2_X1 _4285_ (.A(\fir.p0[8] ),
    .B(\fir.p0[6] ),
    .Z(_3541_));
 XNOR2_X1 _4286_ (.A(_3540_),
    .B(_3541_),
    .ZN(_3542_));
 XNOR2_X1 _4287_ (.A(\fir.p0[4] ),
    .B(_3542_),
    .ZN(_3543_));
 XOR2_X1 _4288_ (.A(_3539_),
    .B(_3543_),
    .Z(_3544_));
 OR2_X1 _4289_ (.A1(\fir.p1[8] ),
    .A2(\fir.p1[7] ),
    .ZN(_3545_));
 NAND2_X1 _4290_ (.A1(\fir.p1[8] ),
    .A2(\fir.p1[7] ),
    .ZN(_3546_));
 AOI22_X1 _4291_ (.A1(\fir.p1[7] ),
    .A2(\fir.p1[6] ),
    .B1(_3545_),
    .B2(_3546_),
    .ZN(_3547_));
 NOR2_X1 _4292_ (.A1(\fir.p1[8] ),
    .A2(_3375_),
    .ZN(_3548_));
 NOR2_X1 _4293_ (.A1(_3547_),
    .A2(_3548_),
    .ZN(_3549_));
 XNOR2_X1 _4294_ (.A(_3544_),
    .B(_3549_),
    .ZN(_3550_));
 XOR2_X1 _4295_ (.A(_3537_),
    .B(_3550_),
    .Z(_3551_));
 XNOR2_X1 _4296_ (.A(_0002_),
    .B(_3377_),
    .ZN(_3552_));
 XNOR2_X1 _4297_ (.A(_3551_),
    .B(_3552_),
    .ZN(_3553_));
 XOR2_X1 _4298_ (.A(_3535_),
    .B(_3553_),
    .Z(_3554_));
 XNOR2_X1 _4299_ (.A(_3533_),
    .B(_3554_),
    .ZN(_3555_));
 XOR2_X1 _4300_ (.A(_3532_),
    .B(_3555_),
    .Z(_3556_));
 XNOR2_X1 _4301_ (.A(_3530_),
    .B(_3556_),
    .ZN(_3557_));
 XNOR2_X1 _4302_ (.A(_3529_),
    .B(_3557_),
    .ZN(_3558_));
 XNOR2_X1 _4303_ (.A(\fir.p2[5] ),
    .B(_3558_),
    .ZN(_3559_));
 XOR2_X1 _4304_ (.A(_3526_),
    .B(_3559_),
    .Z(_3560_));
 XOR2_X1 _4305_ (.A(\fir.p2[7] ),
    .B(\fir.p2[3] ),
    .Z(_3561_));
 XNOR2_X1 _4306_ (.A(_3560_),
    .B(_3561_),
    .ZN(_3562_));
 XOR2_X1 _4307_ (.A(_3525_),
    .B(_3562_),
    .Z(_3563_));
 NAND2_X1 _4308_ (.A1(\fir.p2[6] ),
    .A2(\fir.p2[2] ),
    .ZN(_3564_));
 XOR2_X1 _4309_ (.A(_0008_),
    .B(_3564_),
    .Z(_3565_));
 XNOR2_X1 _4310_ (.A(_3563_),
    .B(_3565_),
    .ZN(_3566_));
 XOR2_X1 _4311_ (.A(_3523_),
    .B(_3566_),
    .Z(_3567_));
 XOR2_X1 _4312_ (.A(_3521_),
    .B(_3567_),
    .Z(_3568_));
 XOR2_X1 _4313_ (.A(_3520_),
    .B(_3568_),
    .Z(_3569_));
 XNOR2_X1 _4314_ (.A(_3518_),
    .B(_3569_),
    .ZN(_3570_));
 XNOR2_X1 _4315_ (.A(_3517_),
    .B(_3570_),
    .ZN(_3571_));
 XOR2_X1 _4316_ (.A(_3516_),
    .B(_3571_),
    .Z(_3572_));
 XOR2_X1 _4317_ (.A(\fir.p4[6] ),
    .B(\fir.p4[5] ),
    .Z(_3573_));
 XNOR2_X1 _4318_ (.A(\fir.p4[4] ),
    .B(_3573_),
    .ZN(_3574_));
 INV_X1 _4319_ (.A(_3574_),
    .ZN(_3575_));
 XNOR2_X1 _4320_ (.A(_3572_),
    .B(_3575_),
    .ZN(_3576_));
 XOR2_X1 _4321_ (.A(_3515_),
    .B(_3576_),
    .Z(_3577_));
 AND2_X1 _4322_ (.A1(\fir.p4[5] ),
    .A2(\fir.p4[4] ),
    .ZN(_3578_));
 AOI21_X1 _4323_ (.A(_3578_),
    .B1(_3403_),
    .B2(\fir.p4[3] ),
    .ZN(_3579_));
 XNOR2_X1 _4324_ (.A(_3200_),
    .B(_3579_),
    .ZN(_3580_));
 XOR2_X1 _4325_ (.A(_3139_),
    .B(_3580_),
    .Z(_3581_));
 XNOR2_X1 _4326_ (.A(_3577_),
    .B(_3581_),
    .ZN(_3582_));
 XOR2_X1 _4327_ (.A(_3513_),
    .B(_3582_),
    .Z(_3583_));
 INV_X1 _4328_ (.A(_3419_),
    .ZN(_3584_));
 NAND2_X1 _4329_ (.A1(\fir.p3[7] ),
    .A2(_3584_),
    .ZN(_3585_));
 XOR2_X1 _4330_ (.A(\fir.p3[6] ),
    .B(\fir.p3[5] ),
    .Z(_3586_));
 XNOR2_X1 _4331_ (.A(\fir.p3[4] ),
    .B(_3586_),
    .ZN(_3587_));
 XOR2_X1 _4332_ (.A(\fir.p3[8] ),
    .B(_3587_),
    .Z(_3588_));
 NOR2_X1 _4333_ (.A1(_3141_),
    .A2(_3409_),
    .ZN(_3589_));
 NOR2_X1 _4334_ (.A1(_3229_),
    .A2(_3410_),
    .ZN(_3590_));
 NOR2_X1 _4335_ (.A1(_3589_),
    .A2(_3590_),
    .ZN(_3591_));
 XNOR2_X1 _4336_ (.A(_3588_),
    .B(_3591_),
    .ZN(_3592_));
 XOR2_X1 _4337_ (.A(_3585_),
    .B(_3592_),
    .Z(_3593_));
 XNOR2_X1 _4338_ (.A(_3583_),
    .B(_3593_),
    .ZN(_3594_));
 XOR2_X1 _4339_ (.A(_3511_),
    .B(_3594_),
    .Z(_3595_));
 AND2_X1 _4340_ (.A1(_3426_),
    .A2(_3431_),
    .ZN(_3596_));
 OAI21_X1 _4341_ (.A(_3327_),
    .B1(\fir.p3[0] ),
    .B2(\fir.p3[2] ),
    .ZN(_3597_));
 AND2_X1 _4342_ (.A1(\fir.p3[5] ),
    .A2(\fir.p3[4] ),
    .ZN(_3598_));
 AOI21_X1 _4343_ (.A(_3598_),
    .B1(_3418_),
    .B2(\fir.p3[3] ),
    .ZN(_3599_));
 XNOR2_X1 _4344_ (.A(_3212_),
    .B(_3599_),
    .ZN(_3600_));
 XNOR2_X1 _4345_ (.A(_3597_),
    .B(_3600_),
    .ZN(_3601_));
 OR2_X1 _4346_ (.A1(_3427_),
    .A2(_3430_),
    .ZN(_3602_));
 OR2_X1 _4347_ (.A1(_3208_),
    .A2(_3429_),
    .ZN(_3603_));
 AOI21_X1 _4348_ (.A(_3601_),
    .B1(_3602_),
    .B2(_3603_),
    .ZN(_3604_));
 AND3_X1 _4349_ (.A1(_3603_),
    .A2(_3602_),
    .A3(_3601_),
    .ZN(_3605_));
 NOR2_X1 _4350_ (.A1(_3604_),
    .A2(_3605_),
    .ZN(_3606_));
 NOR2_X1 _4351_ (.A1(_3415_),
    .A2(_3421_),
    .ZN(_3607_));
 NOR3_X1 _4352_ (.A1(_3416_),
    .A2(_3311_),
    .A3(_3420_),
    .ZN(_3608_));
 OAI21_X1 _4353_ (.A(_3606_),
    .B1(_3607_),
    .B2(_3608_),
    .ZN(_3609_));
 INV_X1 _4354_ (.A(_3609_),
    .ZN(_3610_));
 NOR3_X1 _4355_ (.A1(_3608_),
    .A2(_3607_),
    .A3(_3606_),
    .ZN(_3611_));
 NOR2_X1 _4356_ (.A1(_3610_),
    .A2(_3611_),
    .ZN(_3612_));
 XOR2_X1 _4357_ (.A(_3596_),
    .B(_3612_),
    .Z(_3613_));
 XNOR2_X1 _4358_ (.A(_3595_),
    .B(_3613_),
    .ZN(_3614_));
 XOR2_X1 _4359_ (.A(_3509_),
    .B(_3614_),
    .Z(_3615_));
 OAI21_X1 _4360_ (.A(_3436_),
    .B1(_3438_),
    .B2(_3425_),
    .ZN(_3616_));
 XOR2_X1 _4361_ (.A(_3615_),
    .B(_3616_),
    .Z(_3617_));
 XNOR2_X1 _4362_ (.A(_3507_),
    .B(_3617_),
    .ZN(_3618_));
 XNOR2_X1 _4363_ (.A(_3505_),
    .B(_3618_),
    .ZN(_3619_));
 NAND2_X1 _4364_ (.A1(\fir.p5[7] ),
    .A2(_3619_),
    .ZN(_3620_));
 NOR2_X1 _4365_ (.A1(_3509_),
    .A2(_3614_),
    .ZN(_3621_));
 AOI21_X1 _4366_ (.A(_3621_),
    .B1(_3615_),
    .B2(_3616_),
    .ZN(_3622_));
 NOR2_X1 _4367_ (.A1(_3511_),
    .A2(_3594_),
    .ZN(_3623_));
 AOI21_X1 _4368_ (.A(_3623_),
    .B1(_3595_),
    .B2(_3613_),
    .ZN(_3624_));
 OR2_X1 _4369_ (.A1(_3513_),
    .A2(_3582_),
    .ZN(_3625_));
 NAND2_X1 _4370_ (.A1(_3583_),
    .A2(_3593_),
    .ZN(_3626_));
 NAND2_X1 _4371_ (.A1(_3625_),
    .A2(_3626_),
    .ZN(_3627_));
 OR2_X1 _4372_ (.A1(_3515_),
    .A2(_3576_),
    .ZN(_3628_));
 NAND2_X1 _4373_ (.A1(_3577_),
    .A2(_3581_),
    .ZN(_3629_));
 NAND2_X1 _4374_ (.A1(_3628_),
    .A2(_3629_),
    .ZN(_3630_));
 NOR2_X1 _4375_ (.A1(_3516_),
    .A2(_3571_),
    .ZN(_3631_));
 AND2_X1 _4376_ (.A1(_3572_),
    .A2(_3575_),
    .ZN(_3632_));
 NOR2_X1 _4377_ (.A1(_3631_),
    .A2(_3632_),
    .ZN(_3633_));
 NOR2_X1 _4378_ (.A1(_3517_),
    .A2(_3570_),
    .ZN(_3634_));
 AND2_X1 _4379_ (.A1(_3520_),
    .A2(_3568_),
    .ZN(_3635_));
 AOI21_X1 _4380_ (.A(_3635_),
    .B1(_3569_),
    .B2(_3518_),
    .ZN(_3636_));
 NOR2_X1 _4381_ (.A1(_3523_),
    .A2(_3566_),
    .ZN(_3637_));
 AOI21_X1 _4382_ (.A(_3637_),
    .B1(_3567_),
    .B2(_3521_),
    .ZN(_3638_));
 NOR2_X1 _4383_ (.A1(_0008_),
    .A2(_3564_),
    .ZN(_3639_));
 OR2_X1 _4384_ (.A1(_3525_),
    .A2(_3562_),
    .ZN(_3640_));
 NAND2_X1 _4385_ (.A1(_3563_),
    .A2(_3565_),
    .ZN(_3641_));
 NAND2_X1 _4386_ (.A1(_3640_),
    .A2(_3641_),
    .ZN(_3642_));
 OR2_X1 _4387_ (.A1(_3526_),
    .A2(_3559_),
    .ZN(_3643_));
 NAND2_X1 _4388_ (.A1(_3560_),
    .A2(_3561_),
    .ZN(_3644_));
 NAND2_X1 _4389_ (.A1(_3643_),
    .A2(_3644_),
    .ZN(_3645_));
 NAND2_X1 _4390_ (.A1(\fir.p2[5] ),
    .A2(_3558_),
    .ZN(_3646_));
 NOR2_X1 _4391_ (.A1(_3532_),
    .A2(_3555_),
    .ZN(_3647_));
 NOR2_X1 _4392_ (.A1(_3535_),
    .A2(_3553_),
    .ZN(_3648_));
 AOI21_X1 _4393_ (.A(_3648_),
    .B1(_3554_),
    .B2(_3533_),
    .ZN(_3649_));
 NOR3_X1 _4394_ (.A1(\fir.p1[7] ),
    .A2(_0002_),
    .A3(_3276_),
    .ZN(_3650_));
 NOR2_X1 _4395_ (.A1(_3537_),
    .A2(_3550_),
    .ZN(_3651_));
 AOI21_X1 _4396_ (.A(_3651_),
    .B1(_3551_),
    .B2(_3552_),
    .ZN(_3652_));
 NOR2_X1 _4397_ (.A1(_3539_),
    .A2(_3543_),
    .ZN(_3653_));
 AOI21_X1 _4398_ (.A(_3653_),
    .B1(_3544_),
    .B2(_3549_),
    .ZN(_3654_));
 AND3_X1 _4399_ (.A1(\fir.p0[7] ),
    .A2(\fir.p0[5] ),
    .A3(_3541_),
    .ZN(_3655_));
 AOI21_X1 _4400_ (.A(_3655_),
    .B1(_3542_),
    .B2(\fir.p0[4] ),
    .ZN(_3656_));
 NAND2_X1 _4401_ (.A1(\fir.p0[8] ),
    .A2(\fir.p0[6] ),
    .ZN(_3657_));
 XOR2_X1 _4402_ (.A(\fir.p0[9] ),
    .B(\fir.p0[7] ),
    .Z(_3658_));
 XNOR2_X1 _4403_ (.A(_3657_),
    .B(_3658_),
    .ZN(_3659_));
 XNOR2_X1 _4404_ (.A(\fir.p0[5] ),
    .B(_3659_),
    .ZN(_3660_));
 XOR2_X1 _4405_ (.A(_3656_),
    .B(_3660_),
    .Z(_3661_));
 OR2_X1 _4406_ (.A1(\fir.p1[9] ),
    .A2(\fir.p1[8] ),
    .ZN(_3662_));
 NAND2_X1 _4407_ (.A1(\fir.p1[9] ),
    .A2(\fir.p1[8] ),
    .ZN(_3663_));
 AOI22_X1 _4408_ (.A1(\fir.p1[8] ),
    .A2(\fir.p1[7] ),
    .B1(_3662_),
    .B2(_3663_),
    .ZN(_3664_));
 NOR2_X1 _4409_ (.A1(\fir.p1[9] ),
    .A2(_3546_),
    .ZN(_3665_));
 NOR2_X1 _4410_ (.A1(_3664_),
    .A2(_3665_),
    .ZN(_3666_));
 XNOR2_X1 _4411_ (.A(_3661_),
    .B(_3666_),
    .ZN(_0215_));
 XOR2_X1 _4412_ (.A(_3654_),
    .B(_0215_),
    .Z(_0216_));
 XNOR2_X1 _4413_ (.A(_0001_),
    .B(_3548_),
    .ZN(_0217_));
 XNOR2_X1 _4414_ (.A(_0216_),
    .B(_0217_),
    .ZN(_0218_));
 XOR2_X1 _4415_ (.A(_3652_),
    .B(_0218_),
    .Z(_0219_));
 XNOR2_X1 _4416_ (.A(_3650_),
    .B(_0219_),
    .ZN(_0220_));
 XOR2_X1 _4417_ (.A(_3649_),
    .B(_0220_),
    .Z(_0221_));
 XNOR2_X1 _4418_ (.A(_3647_),
    .B(_0221_),
    .ZN(_0222_));
 AND2_X1 _4419_ (.A1(_3530_),
    .A2(_3556_),
    .ZN(_0223_));
 INV_X1 _4420_ (.A(_3557_),
    .ZN(_0224_));
 AOI21_X1 _4421_ (.A(_0223_),
    .B1(_0224_),
    .B2(_3529_),
    .ZN(_0225_));
 XNOR2_X1 _4422_ (.A(_0222_),
    .B(_0225_),
    .ZN(_0226_));
 XOR2_X1 _4423_ (.A(\fir.p2[6] ),
    .B(_0226_),
    .Z(_0227_));
 XOR2_X1 _4424_ (.A(_3646_),
    .B(_0227_),
    .Z(_0228_));
 XOR2_X1 _4425_ (.A(\fir.p2[8] ),
    .B(\fir.p2[4] ),
    .Z(_0229_));
 XNOR2_X1 _4426_ (.A(_0228_),
    .B(_0229_),
    .ZN(_0230_));
 XNOR2_X1 _4427_ (.A(_3645_),
    .B(_0230_),
    .ZN(_0231_));
 NAND2_X1 _4428_ (.A1(\fir.p2[7] ),
    .A2(\fir.p2[3] ),
    .ZN(_0232_));
 XOR2_X1 _4429_ (.A(_0007_),
    .B(_0232_),
    .Z(_0233_));
 XNOR2_X1 _4430_ (.A(_0231_),
    .B(_0233_),
    .ZN(_0234_));
 XNOR2_X1 _4431_ (.A(_3642_),
    .B(_0234_),
    .ZN(_0235_));
 XNOR2_X1 _4432_ (.A(_3639_),
    .B(_0235_),
    .ZN(_0236_));
 XNOR2_X1 _4433_ (.A(_3638_),
    .B(_0236_),
    .ZN(_0237_));
 XOR2_X1 _4434_ (.A(_3636_),
    .B(_0237_),
    .Z(_0238_));
 XOR2_X1 _4435_ (.A(\fir.p4[9] ),
    .B(_0238_),
    .Z(_0239_));
 XNOR2_X1 _4436_ (.A(_3634_),
    .B(_0239_),
    .ZN(_0240_));
 XOR2_X1 _4437_ (.A(\fir.p4[7] ),
    .B(\fir.p4[6] ),
    .Z(_0241_));
 XNOR2_X1 _4438_ (.A(\fir.p4[5] ),
    .B(_0241_),
    .ZN(_0242_));
 XOR2_X1 _4439_ (.A(_0240_),
    .B(_0242_),
    .Z(_0243_));
 XNOR2_X1 _4440_ (.A(_3633_),
    .B(_0243_),
    .ZN(_0244_));
 AND2_X1 _4441_ (.A1(\fir.p4[6] ),
    .A2(\fir.p4[5] ),
    .ZN(_0245_));
 AOI21_X1 _4442_ (.A(_0245_),
    .B1(_3573_),
    .B2(\fir.p4[4] ),
    .ZN(_0246_));
 XNOR2_X1 _4443_ (.A(_3307_),
    .B(_0246_),
    .ZN(_0247_));
 XOR2_X1 _4444_ (.A(_3311_),
    .B(_0247_),
    .Z(_0248_));
 XNOR2_X1 _4445_ (.A(_0244_),
    .B(_0248_),
    .ZN(_0249_));
 XNOR2_X1 _4446_ (.A(_3630_),
    .B(_0249_),
    .ZN(_0250_));
 INV_X1 _4447_ (.A(_3587_),
    .ZN(_0251_));
 NAND2_X1 _4448_ (.A1(\fir.p3[8] ),
    .A2(_0251_),
    .ZN(_0252_));
 XOR2_X1 _4449_ (.A(\fir.p3[7] ),
    .B(\fir.p3[6] ),
    .Z(_0253_));
 XNOR2_X1 _4450_ (.A(\fir.p3[5] ),
    .B(_0253_),
    .ZN(_0254_));
 XOR2_X1 _4451_ (.A(\fir.p3[9] ),
    .B(_0254_),
    .Z(_0255_));
 NOR2_X1 _4452_ (.A1(_3200_),
    .A2(_3579_),
    .ZN(_0256_));
 NOR2_X1 _4453_ (.A1(_3139_),
    .A2(_3580_),
    .ZN(_0257_));
 NOR2_X1 _4454_ (.A1(_0256_),
    .A2(_0257_),
    .ZN(_0258_));
 XNOR2_X1 _4455_ (.A(_0255_),
    .B(_0258_),
    .ZN(_0259_));
 XOR2_X1 _4456_ (.A(_0252_),
    .B(_0259_),
    .Z(_0260_));
 XNOR2_X1 _4457_ (.A(_0250_),
    .B(_0260_),
    .ZN(_0261_));
 XNOR2_X1 _4458_ (.A(_3627_),
    .B(_0261_),
    .ZN(_0262_));
 NOR2_X1 _4459_ (.A1(_3212_),
    .A2(_3599_),
    .ZN(_0263_));
 NOR2_X1 _4460_ (.A1(_3597_),
    .A2(_3600_),
    .ZN(_0264_));
 NOR2_X1 _4461_ (.A1(_0263_),
    .A2(_0264_),
    .ZN(_0265_));
 AND2_X1 _4462_ (.A1(\fir.p3[6] ),
    .A2(\fir.p3[5] ),
    .ZN(_0266_));
 AOI21_X1 _4463_ (.A(_0266_),
    .B1(_3586_),
    .B2(\fir.p3[4] ),
    .ZN(_0267_));
 XNOR2_X1 _4464_ (.A(_3318_),
    .B(_0267_),
    .ZN(_0268_));
 XOR2_X1 _4465_ (.A(_3330_),
    .B(_0268_),
    .Z(_0269_));
 XNOR2_X1 _4466_ (.A(_0265_),
    .B(_0269_),
    .ZN(_0270_));
 NOR2_X1 _4467_ (.A1(_3585_),
    .A2(_3592_),
    .ZN(_0271_));
 NOR2_X1 _4468_ (.A1(_3588_),
    .A2(_3591_),
    .ZN(_0272_));
 OAI21_X1 _4469_ (.A(_0270_),
    .B1(_0271_),
    .B2(_0272_),
    .ZN(_0273_));
 OR3_X1 _4470_ (.A1(_0272_),
    .A2(_0271_),
    .A3(_0270_),
    .ZN(_0274_));
 AND2_X1 _4471_ (.A1(_0273_),
    .A2(_0274_),
    .ZN(_0275_));
 XOR2_X1 _4472_ (.A(_3604_),
    .B(_0275_),
    .Z(_0276_));
 XNOR2_X1 _4473_ (.A(_0262_),
    .B(_0276_),
    .ZN(_0277_));
 XOR2_X1 _4474_ (.A(_3624_),
    .B(_0277_),
    .Z(_0278_));
 AOI21_X1 _4475_ (.A(_3610_),
    .B1(_3612_),
    .B2(_3596_),
    .ZN(_0279_));
 XNOR2_X1 _4476_ (.A(_0278_),
    .B(_0279_),
    .ZN(_0280_));
 XNOR2_X1 _4477_ (.A(_3622_),
    .B(_0280_),
    .ZN(_0281_));
 INV_X1 _4478_ (.A(_3507_),
    .ZN(_0282_));
 AND2_X1 _4479_ (.A1(_0282_),
    .A2(_3617_),
    .ZN(_0283_));
 OR2_X1 _4480_ (.A1(_3338_),
    .A2(_3442_),
    .ZN(_0284_));
 NOR2_X1 _4481_ (.A1(_3468_),
    .A2(_3502_),
    .ZN(_0285_));
 AND2_X1 _4482_ (.A1(_3338_),
    .A2(_3442_),
    .ZN(_0286_));
 OAI21_X1 _4483_ (.A(_0284_),
    .B1(_0285_),
    .B2(_0286_),
    .ZN(_0287_));
 AOI21_X1 _4484_ (.A(_0283_),
    .B1(_3618_),
    .B2(_0287_),
    .ZN(_0288_));
 XNOR2_X1 _4485_ (.A(_0281_),
    .B(_0288_),
    .ZN(_0289_));
 XNOR2_X1 _4486_ (.A(\fir.p5[8] ),
    .B(_0289_),
    .ZN(_0290_));
 NOR2_X1 _4487_ (.A1(_3620_),
    .A2(_0290_),
    .ZN(_0291_));
 XOR2_X1 _4488_ (.A(_3620_),
    .B(_0290_),
    .Z(_0292_));
 XOR2_X1 _4489_ (.A(\fir.p5[6] ),
    .B(\fir.p5[4] ),
    .Z(_0293_));
 AOI21_X1 _4490_ (.A(_0291_),
    .B1(_0292_),
    .B2(_0293_),
    .ZN(_0294_));
 XOR2_X1 _4491_ (.A(\fir.p5[7] ),
    .B(\fir.p5[5] ),
    .Z(_0295_));
 NAND2_X1 _4492_ (.A1(\fir.p5[8] ),
    .A2(_0289_),
    .ZN(_0296_));
 XNOR2_X1 _4493_ (.A(_0282_),
    .B(_3617_),
    .ZN(_0297_));
 INV_X1 _4494_ (.A(_0279_),
    .ZN(_0298_));
 XNOR2_X1 _4495_ (.A(_0278_),
    .B(_0298_),
    .ZN(_0299_));
 OAI22_X1 _4496_ (.A1(_3505_),
    .A2(_0297_),
    .B1(_3622_),
    .B2(_0299_),
    .ZN(_0300_));
 NAND2_X1 _4497_ (.A1(_3622_),
    .A2(_0299_),
    .ZN(_0301_));
 AOI22_X1 _4498_ (.A1(_0283_),
    .A2(_0281_),
    .B1(_0300_),
    .B2(_0301_),
    .ZN(_0302_));
 NOR2_X1 _4499_ (.A1(_3624_),
    .A2(_0277_),
    .ZN(_0303_));
 AOI21_X1 _4500_ (.A(_0303_),
    .B1(_0278_),
    .B2(_0298_),
    .ZN(_0304_));
 NAND2_X1 _4501_ (.A1(_3604_),
    .A2(_0275_),
    .ZN(_0305_));
 NAND2_X1 _4502_ (.A1(_0273_),
    .A2(_0305_),
    .ZN(_0306_));
 AOI21_X1 _4503_ (.A(_0261_),
    .B1(_3626_),
    .B2(_3625_),
    .ZN(_0307_));
 AOI21_X1 _4504_ (.A(_0307_),
    .B1(_0262_),
    .B2(_0276_),
    .ZN(_0308_));
 OAI21_X1 _4505_ (.A(_0269_),
    .B1(_0264_),
    .B2(_0263_),
    .ZN(_0309_));
 NOR2_X1 _4506_ (.A1(_3318_),
    .A2(_0267_),
    .ZN(_0310_));
 NOR2_X1 _4507_ (.A1(_3330_),
    .A2(_0268_),
    .ZN(_0311_));
 NOR2_X1 _4508_ (.A1(_0310_),
    .A2(_0311_),
    .ZN(_0312_));
 AND2_X1 _4509_ (.A1(\fir.p3[7] ),
    .A2(\fir.p3[6] ),
    .ZN(_0313_));
 AOI21_X1 _4510_ (.A(_0313_),
    .B1(_0253_),
    .B2(\fir.p3[5] ),
    .ZN(_0314_));
 XNOR2_X1 _4511_ (.A(_3419_),
    .B(_0314_),
    .ZN(_0315_));
 XOR2_X1 _4512_ (.A(_3429_),
    .B(_0315_),
    .Z(_0316_));
 XNOR2_X1 _4513_ (.A(_0312_),
    .B(_0316_),
    .ZN(_0317_));
 NOR2_X1 _4514_ (.A1(_0255_),
    .A2(_0258_),
    .ZN(_0318_));
 NOR2_X1 _4515_ (.A1(_0252_),
    .A2(_0259_),
    .ZN(_0319_));
 NOR2_X1 _4516_ (.A1(_0318_),
    .A2(_0319_),
    .ZN(_0320_));
 XNOR2_X1 _4517_ (.A(_0317_),
    .B(_0320_),
    .ZN(_0321_));
 XNOR2_X1 _4518_ (.A(_0309_),
    .B(_0321_),
    .ZN(_0322_));
 AOI21_X1 _4519_ (.A(_0249_),
    .B1(_3629_),
    .B2(_3628_),
    .ZN(_0323_));
 AOI21_X1 _4520_ (.A(_0323_),
    .B1(_0250_),
    .B2(_0260_),
    .ZN(_0324_));
 INV_X1 _4521_ (.A(_0254_),
    .ZN(_0325_));
 NAND2_X1 _4522_ (.A1(\fir.p3[9] ),
    .A2(_0325_),
    .ZN(_0326_));
 XOR2_X1 _4523_ (.A(\fir.p3[8] ),
    .B(\fir.p3[7] ),
    .Z(_0327_));
 XNOR2_X1 _4524_ (.A(\fir.p3[6] ),
    .B(_0327_),
    .ZN(_0328_));
 XOR2_X1 _4525_ (.A(\fir.p3[10] ),
    .B(_0328_),
    .Z(_0329_));
 NOR2_X1 _4526_ (.A1(_3307_),
    .A2(_0246_),
    .ZN(_0330_));
 NOR2_X1 _4527_ (.A1(_3311_),
    .A2(_0247_),
    .ZN(_0331_));
 NOR2_X1 _4528_ (.A1(_0330_),
    .A2(_0331_),
    .ZN(_0332_));
 XNOR2_X1 _4529_ (.A(_0329_),
    .B(_0332_),
    .ZN(_0333_));
 XOR2_X1 _4530_ (.A(_0326_),
    .B(_0333_),
    .Z(_0334_));
 OAI21_X1 _4531_ (.A(_0243_),
    .B1(_3632_),
    .B2(_3631_),
    .ZN(_0335_));
 INV_X1 _4532_ (.A(_0335_),
    .ZN(_0336_));
 AOI21_X1 _4533_ (.A(_0336_),
    .B1(_0244_),
    .B2(_0248_),
    .ZN(_0337_));
 AND2_X1 _4534_ (.A1(\fir.p4[7] ),
    .A2(\fir.p4[6] ),
    .ZN(_0338_));
 AOI21_X1 _4535_ (.A(_0338_),
    .B1(_0241_),
    .B2(\fir.p4[5] ),
    .ZN(_0339_));
 XNOR2_X1 _4536_ (.A(_3404_),
    .B(_0339_),
    .ZN(_0340_));
 XOR2_X1 _4537_ (.A(_3409_),
    .B(_0340_),
    .Z(_0341_));
 INV_X1 _4538_ (.A(_0341_),
    .ZN(_0342_));
 NAND2_X1 _4539_ (.A1(_3634_),
    .A2(_0239_),
    .ZN(_0343_));
 OAI21_X1 _4540_ (.A(_0343_),
    .B1(_0240_),
    .B2(_0242_),
    .ZN(_0344_));
 XOR2_X1 _4541_ (.A(\fir.p4[8] ),
    .B(\fir.p4[7] ),
    .Z(_0345_));
 XNOR2_X1 _4542_ (.A(\fir.p4[6] ),
    .B(_0345_),
    .ZN(_0346_));
 NAND2_X1 _4543_ (.A1(\fir.p4[9] ),
    .A2(_0238_),
    .ZN(_0347_));
 AOI21_X1 _4544_ (.A(_0234_),
    .B1(_3641_),
    .B2(_3640_),
    .ZN(_0348_));
 AOI21_X1 _4545_ (.A(_0348_),
    .B1(_0235_),
    .B2(_3639_),
    .ZN(_0349_));
 NOR2_X1 _4546_ (.A1(_0007_),
    .A2(_0232_),
    .ZN(_0350_));
 AOI21_X1 _4547_ (.A(_0230_),
    .B1(_3644_),
    .B2(_3643_),
    .ZN(_0351_));
 AOI21_X1 _4548_ (.A(_0351_),
    .B1(_0231_),
    .B2(_0233_),
    .ZN(_0352_));
 NAND2_X1 _4549_ (.A1(\fir.p2[8] ),
    .A2(\fir.p2[4] ),
    .ZN(_0353_));
 XOR2_X1 _4550_ (.A(_0006_),
    .B(_0353_),
    .Z(_0354_));
 NOR2_X1 _4551_ (.A1(_3646_),
    .A2(_0227_),
    .ZN(_0355_));
 AOI21_X1 _4552_ (.A(_0355_),
    .B1(_0228_),
    .B2(_0229_),
    .ZN(_0356_));
 XNOR2_X1 _4553_ (.A(\fir.p2[9] ),
    .B(\fir.p2[5] ),
    .ZN(_0357_));
 OR2_X1 _4554_ (.A1(_0005_),
    .A2(_0226_),
    .ZN(_0358_));
 NAND2_X1 _4555_ (.A1(_3647_),
    .A2(_0221_),
    .ZN(_0359_));
 NAND2_X1 _4556_ (.A1(_3530_),
    .A2(_3556_),
    .ZN(_0360_));
 OAI21_X1 _4557_ (.A(_0359_),
    .B1(_0222_),
    .B2(_0360_),
    .ZN(_0361_));
 NOR2_X1 _4558_ (.A1(_3557_),
    .A2(_0222_),
    .ZN(_0362_));
 AOI21_X1 _4559_ (.A(_0361_),
    .B1(_0362_),
    .B2(_3529_),
    .ZN(_0363_));
 NOR2_X1 _4560_ (.A1(_3649_),
    .A2(_0220_),
    .ZN(_0364_));
 NOR2_X1 _4561_ (.A1(_3652_),
    .A2(_0218_),
    .ZN(_0365_));
 AOI21_X1 _4562_ (.A(_0365_),
    .B1(_0219_),
    .B2(_3650_),
    .ZN(_0366_));
 NOR3_X1 _4563_ (.A1(\fir.p1[8] ),
    .A2(_0001_),
    .A3(_3375_),
    .ZN(_0367_));
 NOR2_X1 _4564_ (.A1(_3654_),
    .A2(_0215_),
    .ZN(_0368_));
 AOI21_X1 _4565_ (.A(_0368_),
    .B1(_0216_),
    .B2(_0217_),
    .ZN(_0369_));
 XNOR2_X1 _4566_ (.A(_0000_),
    .B(_3665_),
    .ZN(_0370_));
 NOR2_X1 _4567_ (.A1(_3656_),
    .A2(_3660_),
    .ZN(_0371_));
 AOI21_X1 _4568_ (.A(_0371_),
    .B1(_3661_),
    .B2(_3666_),
    .ZN(_0372_));
 OR2_X1 _4569_ (.A1(\fir.p1[9] ),
    .A2(\fir.p1[10] ),
    .ZN(_0373_));
 NAND2_X1 _4570_ (.A1(\fir.p1[9] ),
    .A2(\fir.p1[10] ),
    .ZN(_0374_));
 AOI22_X1 _4571_ (.A1(\fir.p1[9] ),
    .A2(\fir.p1[8] ),
    .B1(_0373_),
    .B2(_0374_),
    .ZN(_0375_));
 NOR2_X1 _4572_ (.A1(\fir.p1[10] ),
    .A2(_3663_),
    .ZN(_0376_));
 NOR2_X1 _4573_ (.A1(_0375_),
    .A2(_0376_),
    .ZN(_0377_));
 NAND2_X1 _4574_ (.A1(\fir.p0[9] ),
    .A2(\fir.p0[7] ),
    .ZN(_0378_));
 XOR2_X1 _4575_ (.A(\fir.p0[8] ),
    .B(\fir.p0[10] ),
    .Z(_0379_));
 XNOR2_X1 _4576_ (.A(_0378_),
    .B(_0379_),
    .ZN(_0380_));
 XNOR2_X1 _4577_ (.A(\fir.p0[6] ),
    .B(_0380_),
    .ZN(_0381_));
 NAND2_X1 _4578_ (.A1(\fir.p0[5] ),
    .A2(_3659_),
    .ZN(_0382_));
 NAND3_X1 _4579_ (.A1(\fir.p0[8] ),
    .A2(\fir.p0[6] ),
    .A3(_3658_),
    .ZN(_0383_));
 AOI21_X1 _4580_ (.A(_0381_),
    .B1(_0382_),
    .B2(_0383_),
    .ZN(_0384_));
 AND3_X1 _4581_ (.A1(_0383_),
    .A2(_0382_),
    .A3(_0381_),
    .ZN(_0385_));
 NOR2_X1 _4582_ (.A1(_0384_),
    .A2(_0385_),
    .ZN(_0386_));
 XNOR2_X1 _4583_ (.A(_0377_),
    .B(_0386_),
    .ZN(_0387_));
 XOR2_X1 _4584_ (.A(_0372_),
    .B(_0387_),
    .Z(_0388_));
 XNOR2_X1 _4585_ (.A(_0370_),
    .B(_0388_),
    .ZN(_0389_));
 XOR2_X1 _4586_ (.A(_0369_),
    .B(_0389_),
    .Z(_0390_));
 XNOR2_X1 _4587_ (.A(_0367_),
    .B(_0390_),
    .ZN(_0391_));
 XOR2_X1 _4588_ (.A(_0366_),
    .B(_0391_),
    .Z(_0392_));
 XNOR2_X1 _4589_ (.A(_0364_),
    .B(_0392_),
    .ZN(_0393_));
 XNOR2_X1 _4590_ (.A(_0363_),
    .B(_0393_),
    .ZN(_0394_));
 XOR2_X1 _4591_ (.A(\fir.p2[7] ),
    .B(_0394_),
    .Z(_0395_));
 XOR2_X1 _4592_ (.A(_0358_),
    .B(_0395_),
    .Z(_0396_));
 XNOR2_X1 _4593_ (.A(_0357_),
    .B(_0396_),
    .ZN(_0397_));
 XNOR2_X1 _4594_ (.A(_0356_),
    .B(_0397_),
    .ZN(_0398_));
 XNOR2_X1 _4595_ (.A(_0354_),
    .B(_0398_),
    .ZN(_0399_));
 XOR2_X1 _4596_ (.A(_0352_),
    .B(_0399_),
    .Z(_0400_));
 XNOR2_X1 _4597_ (.A(_0350_),
    .B(_0400_),
    .ZN(_0401_));
 XNOR2_X1 _4598_ (.A(_0349_),
    .B(_0401_),
    .ZN(_0402_));
 OR2_X1 _4599_ (.A1(_3638_),
    .A2(_0236_),
    .ZN(_0403_));
 OAI21_X1 _4600_ (.A(_0403_),
    .B1(_0237_),
    .B2(_3636_),
    .ZN(_0404_));
 XNOR2_X1 _4601_ (.A(_0402_),
    .B(_0404_),
    .ZN(_0405_));
 XOR2_X1 _4602_ (.A(\fir.p4[10] ),
    .B(_0405_),
    .Z(_0406_));
 XNOR2_X1 _4603_ (.A(_0347_),
    .B(_0406_),
    .ZN(_0407_));
 XNOR2_X1 _4604_ (.A(_0346_),
    .B(_0407_),
    .ZN(_0408_));
 XNOR2_X1 _4605_ (.A(_0344_),
    .B(_0408_),
    .ZN(_0409_));
 XNOR2_X1 _4606_ (.A(_0342_),
    .B(_0409_),
    .ZN(_0410_));
 XOR2_X1 _4607_ (.A(_0337_),
    .B(_0410_),
    .Z(_0411_));
 XNOR2_X1 _4608_ (.A(_0334_),
    .B(_0411_),
    .ZN(_0412_));
 XOR2_X1 _4609_ (.A(_0324_),
    .B(_0412_),
    .Z(_0413_));
 XNOR2_X1 _4610_ (.A(_0322_),
    .B(_0413_),
    .ZN(_0414_));
 XOR2_X1 _4611_ (.A(_0308_),
    .B(_0414_),
    .Z(_0415_));
 XNOR2_X1 _4612_ (.A(_0306_),
    .B(_0415_),
    .ZN(_0416_));
 XOR2_X1 _4613_ (.A(_0304_),
    .B(_0416_),
    .Z(_0417_));
 XNOR2_X1 _4614_ (.A(_0302_),
    .B(_0417_),
    .ZN(_0418_));
 XNOR2_X1 _4615_ (.A(\fir.p5[9] ),
    .B(_0418_),
    .ZN(_0419_));
 XOR2_X1 _4616_ (.A(_0296_),
    .B(_0419_),
    .Z(_0420_));
 XNOR2_X1 _4617_ (.A(_0295_),
    .B(_0420_),
    .ZN(_0421_));
 NOR2_X1 _4618_ (.A1(_0294_),
    .A2(_0421_),
    .ZN(_0422_));
 NAND2_X1 _4619_ (.A1(\fir.p5[6] ),
    .A2(\fir.p5[4] ),
    .ZN(_0423_));
 XOR2_X1 _4620_ (.A(_0012_),
    .B(_0423_),
    .Z(_0424_));
 XOR2_X1 _4621_ (.A(_0294_),
    .B(_0421_),
    .Z(_0425_));
 AOI21_X1 _4622_ (.A(_0422_),
    .B1(_0424_),
    .B2(_0425_),
    .ZN(_0426_));
 NAND2_X1 _4623_ (.A1(\fir.p5[7] ),
    .A2(\fir.p5[5] ),
    .ZN(_0427_));
 XOR2_X1 _4624_ (.A(_0022_),
    .B(_0427_),
    .Z(_0428_));
 NOR2_X1 _4625_ (.A1(_0296_),
    .A2(_0419_),
    .ZN(_0429_));
 AOI21_X1 _4626_ (.A(_0429_),
    .B1(_0420_),
    .B2(_0295_),
    .ZN(_0430_));
 XOR2_X1 _4627_ (.A(\fir.p5[8] ),
    .B(\fir.p5[6] ),
    .Z(_0431_));
 INV_X1 _4628_ (.A(_0021_),
    .ZN(_0432_));
 NAND2_X1 _4629_ (.A1(_0432_),
    .A2(_0418_),
    .ZN(_0433_));
 INV_X1 _4630_ (.A(net229),
    .ZN(_0434_));
 OR2_X1 _4631_ (.A1(_0304_),
    .A2(_0416_),
    .ZN(_0435_));
 AND2_X1 _4632_ (.A1(_0304_),
    .A2(_0416_),
    .ZN(_0436_));
 OAI21_X1 _4633_ (.A(_0435_),
    .B1(_0436_),
    .B2(_0302_),
    .ZN(_0437_));
 NOR2_X1 _4634_ (.A1(_0308_),
    .A2(_0414_),
    .ZN(_0438_));
 AOI21_X1 _4635_ (.A(_0438_),
    .B1(_0415_),
    .B2(_0306_),
    .ZN(_0439_));
 OAI21_X1 _4636_ (.A(_0317_),
    .B1(_0319_),
    .B2(_0318_),
    .ZN(_0440_));
 INV_X1 _4637_ (.A(_0321_),
    .ZN(_0441_));
 OAI21_X1 _4638_ (.A(_0440_),
    .B1(_0441_),
    .B2(_0309_),
    .ZN(_0442_));
 NOR2_X1 _4639_ (.A1(_0324_),
    .A2(_0412_),
    .ZN(_0443_));
 AOI21_X1 _4640_ (.A(_0443_),
    .B1(_0413_),
    .B2(_0322_),
    .ZN(_0444_));
 INV_X1 _4641_ (.A(_0316_),
    .ZN(_0445_));
 NOR2_X1 _4642_ (.A1(_0312_),
    .A2(_0445_),
    .ZN(_0446_));
 NOR2_X1 _4643_ (.A1(_3419_),
    .A2(_0314_),
    .ZN(_0447_));
 NOR2_X1 _4644_ (.A1(_3429_),
    .A2(_0315_),
    .ZN(_0448_));
 NOR2_X1 _4645_ (.A1(_0447_),
    .A2(_0448_),
    .ZN(_0449_));
 AND2_X1 _4646_ (.A1(\fir.p3[8] ),
    .A2(\fir.p3[7] ),
    .ZN(_0450_));
 AOI21_X1 _4647_ (.A(_0450_),
    .B1(_0327_),
    .B2(\fir.p3[6] ),
    .ZN(_0451_));
 XNOR2_X1 _4648_ (.A(_3587_),
    .B(_0451_),
    .ZN(_0452_));
 XOR2_X1 _4649_ (.A(_3599_),
    .B(_0452_),
    .Z(_0453_));
 XNOR2_X1 _4650_ (.A(_0449_),
    .B(_0453_),
    .ZN(_0454_));
 NOR2_X1 _4651_ (.A1(_0326_),
    .A2(_0333_),
    .ZN(_0455_));
 NOR2_X1 _4652_ (.A1(_0329_),
    .A2(_0332_),
    .ZN(_0456_));
 OAI21_X1 _4653_ (.A(_0454_),
    .B1(_0455_),
    .B2(_0456_),
    .ZN(_0457_));
 OR3_X1 _4654_ (.A1(_0456_),
    .A2(_0455_),
    .A3(_0454_),
    .ZN(_0458_));
 AND2_X1 _4655_ (.A1(_0457_),
    .A2(_0458_),
    .ZN(_0459_));
 XOR2_X1 _4656_ (.A(_0446_),
    .B(_0459_),
    .Z(_0460_));
 NOR2_X1 _4657_ (.A1(_0337_),
    .A2(_0410_),
    .ZN(_0461_));
 AOI21_X1 _4658_ (.A(_0461_),
    .B1(_0411_),
    .B2(_0334_),
    .ZN(_0462_));
 INV_X1 _4659_ (.A(_0328_),
    .ZN(_0463_));
 NAND2_X1 _4660_ (.A1(\fir.p3[10] ),
    .A2(_0463_),
    .ZN(_0464_));
 INV_X1 _4661_ (.A(net430),
    .ZN(_0465_));
 XOR2_X1 _4662_ (.A(\fir.p3[9] ),
    .B(\fir.p3[8] ),
    .Z(_0466_));
 XNOR2_X1 _4663_ (.A(\fir.p3[7] ),
    .B(_0466_),
    .ZN(_0467_));
 XNOR2_X1 _4664_ (.A(_0465_),
    .B(_0467_),
    .ZN(_0468_));
 NOR2_X1 _4665_ (.A1(_3404_),
    .A2(_0339_),
    .ZN(_0469_));
 NOR2_X1 _4666_ (.A1(_3409_),
    .A2(_0340_),
    .ZN(_0470_));
 NOR2_X1 _4667_ (.A1(_0469_),
    .A2(_0470_),
    .ZN(_0471_));
 XNOR2_X1 _4668_ (.A(_0468_),
    .B(_0471_),
    .ZN(_0472_));
 XOR2_X1 _4669_ (.A(_0464_),
    .B(_0472_),
    .Z(_0473_));
 INV_X1 _4670_ (.A(_0473_),
    .ZN(_0474_));
 NAND2_X1 _4671_ (.A1(_0344_),
    .A2(_0408_),
    .ZN(_0475_));
 OAI21_X1 _4672_ (.A(_0475_),
    .B1(_0409_),
    .B2(_0342_),
    .ZN(_0476_));
 AND2_X1 _4673_ (.A1(\fir.p4[8] ),
    .A2(\fir.p4[7] ),
    .ZN(_0477_));
 AOI21_X1 _4674_ (.A(_0477_),
    .B1(_0345_),
    .B2(\fir.p4[6] ),
    .ZN(_0478_));
 XNOR2_X1 _4675_ (.A(_3574_),
    .B(_0478_),
    .ZN(_0479_));
 XOR2_X1 _4676_ (.A(_3579_),
    .B(_0479_),
    .Z(_0480_));
 INV_X1 _4677_ (.A(_0346_),
    .ZN(_0481_));
 NAND2_X1 _4678_ (.A1(_0481_),
    .A2(_0407_),
    .ZN(_0482_));
 INV_X1 _4679_ (.A(_0406_),
    .ZN(_0483_));
 OAI21_X1 _4680_ (.A(_0482_),
    .B1(_0483_),
    .B2(_0347_),
    .ZN(_0484_));
 XOR2_X1 _4681_ (.A(\fir.p4[9] ),
    .B(\fir.p4[8] ),
    .Z(_0485_));
 XNOR2_X1 _4682_ (.A(\fir.p4[7] ),
    .B(_0485_),
    .ZN(_0486_));
 NAND2_X1 _4683_ (.A1(\fir.p4[10] ),
    .A2(_0405_),
    .ZN(_0487_));
 INV_X1 _4684_ (.A(net444),
    .ZN(_0488_));
 NOR3_X1 _4685_ (.A1(_3636_),
    .A2(_0237_),
    .A3(_0402_),
    .ZN(_0489_));
 OR2_X1 _4686_ (.A1(_0349_),
    .A2(_0401_),
    .ZN(_0490_));
 OAI21_X1 _4687_ (.A(_0490_),
    .B1(_0402_),
    .B2(_0403_),
    .ZN(_0491_));
 OR2_X1 _4688_ (.A1(_0489_),
    .A2(_0491_),
    .ZN(_0492_));
 NOR2_X1 _4689_ (.A1(_0352_),
    .A2(_0399_),
    .ZN(_0493_));
 AOI21_X1 _4690_ (.A(_0493_),
    .B1(_0400_),
    .B2(_0350_),
    .ZN(_0494_));
 NOR2_X1 _4691_ (.A1(_0006_),
    .A2(_0353_),
    .ZN(_0495_));
 INV_X1 _4692_ (.A(_0397_),
    .ZN(_0496_));
 NOR2_X1 _4693_ (.A1(_0356_),
    .A2(_0496_),
    .ZN(_0497_));
 AOI21_X1 _4694_ (.A(_0497_),
    .B1(_0398_),
    .B2(_0354_),
    .ZN(_0498_));
 NAND2_X1 _4695_ (.A1(\fir.p2[9] ),
    .A2(\fir.p2[5] ),
    .ZN(_0499_));
 XOR2_X1 _4696_ (.A(_0019_),
    .B(_0499_),
    .Z(_0500_));
 NOR2_X1 _4697_ (.A1(_0358_),
    .A2(_0395_),
    .ZN(_0501_));
 INV_X1 _4698_ (.A(_0357_),
    .ZN(_0502_));
 AOI21_X1 _4699_ (.A(_0501_),
    .B1(_0396_),
    .B2(_0502_),
    .ZN(_0503_));
 XOR2_X1 _4700_ (.A(\fir.p2[6] ),
    .B(\fir.p2[10] ),
    .Z(_0504_));
 OR2_X1 _4701_ (.A1(_0018_),
    .A2(_0394_),
    .ZN(_0505_));
 NAND2_X1 _4702_ (.A1(_0364_),
    .A2(_0392_),
    .ZN(_0506_));
 OAI21_X1 _4703_ (.A(_0506_),
    .B1(_0393_),
    .B2(_0363_),
    .ZN(_0507_));
 NOR2_X1 _4704_ (.A1(_0366_),
    .A2(_0391_),
    .ZN(_0508_));
 NOR2_X1 _4705_ (.A1(_0369_),
    .A2(_0389_),
    .ZN(_0509_));
 AOI21_X1 _4706_ (.A(_0509_),
    .B1(_0390_),
    .B2(_0367_),
    .ZN(_0510_));
 NOR3_X1 _4707_ (.A1(\fir.p1[9] ),
    .A2(_0000_),
    .A3(_3546_),
    .ZN(_0511_));
 NOR2_X1 _4708_ (.A1(_0372_),
    .A2(_0387_),
    .ZN(_0512_));
 AOI21_X1 _4709_ (.A(_0512_),
    .B1(_0388_),
    .B2(_0370_),
    .ZN(_0513_));
 XNOR2_X1 _4710_ (.A(_0017_),
    .B(_0376_),
    .ZN(_0514_));
 AOI21_X1 _4711_ (.A(_0384_),
    .B1(_0386_),
    .B2(_0377_),
    .ZN(_0515_));
 XNOR2_X1 _4712_ (.A(\fir.p1[11] ),
    .B(\fir.p1[10] ),
    .ZN(_0516_));
 XNOR2_X1 _4713_ (.A(_0374_),
    .B(_0516_),
    .ZN(_0517_));
 NAND2_X1 _4714_ (.A1(\fir.p0[8] ),
    .A2(\fir.p0[10] ),
    .ZN(_0518_));
 XOR2_X1 _4715_ (.A(\fir.p0[9] ),
    .B(\fir.p0[11] ),
    .Z(_0519_));
 XNOR2_X1 _4716_ (.A(_0518_),
    .B(_0519_),
    .ZN(_0520_));
 XNOR2_X1 _4717_ (.A(\fir.p0[7] ),
    .B(_0520_),
    .ZN(_0521_));
 NAND2_X1 _4718_ (.A1(\fir.p0[6] ),
    .A2(_0380_),
    .ZN(_0522_));
 NAND3_X1 _4719_ (.A1(\fir.p0[9] ),
    .A2(\fir.p0[7] ),
    .A3(_0379_),
    .ZN(_0523_));
 AOI21_X1 _4720_ (.A(_0521_),
    .B1(_0522_),
    .B2(_0523_),
    .ZN(_0524_));
 AND3_X1 _4721_ (.A1(_0523_),
    .A2(_0522_),
    .A3(_0521_),
    .ZN(_0525_));
 OR2_X1 _4722_ (.A1(_0524_),
    .A2(_0525_),
    .ZN(_0526_));
 XNOR2_X1 _4723_ (.A(_0517_),
    .B(_0526_),
    .ZN(_0527_));
 XOR2_X1 _4724_ (.A(_0515_),
    .B(_0527_),
    .Z(_0528_));
 XNOR2_X1 _4725_ (.A(_0514_),
    .B(_0528_),
    .ZN(_0529_));
 XOR2_X1 _4726_ (.A(_0513_),
    .B(_0529_),
    .Z(_0530_));
 XNOR2_X1 _4727_ (.A(_0511_),
    .B(_0530_),
    .ZN(_0531_));
 XOR2_X1 _4728_ (.A(_0510_),
    .B(_0531_),
    .Z(_0532_));
 XNOR2_X1 _4729_ (.A(_0508_),
    .B(_0532_),
    .ZN(_0533_));
 XOR2_X1 _4730_ (.A(_0507_),
    .B(_0533_),
    .Z(_0534_));
 XOR2_X1 _4731_ (.A(\fir.p2[8] ),
    .B(_0534_),
    .Z(_0535_));
 XOR2_X1 _4732_ (.A(_0505_),
    .B(_0535_),
    .Z(_0536_));
 XNOR2_X1 _4733_ (.A(_0504_),
    .B(_0536_),
    .ZN(_0537_));
 XOR2_X1 _4734_ (.A(_0503_),
    .B(_0537_),
    .Z(_0538_));
 XNOR2_X1 _4735_ (.A(_0500_),
    .B(_0538_),
    .ZN(_0539_));
 XOR2_X1 _4736_ (.A(_0498_),
    .B(_0539_),
    .Z(_0540_));
 XNOR2_X1 _4737_ (.A(_0495_),
    .B(_0540_),
    .ZN(_0541_));
 XOR2_X1 _4738_ (.A(_0494_),
    .B(_0541_),
    .Z(_0542_));
 XNOR2_X1 _4739_ (.A(_0492_),
    .B(_0542_),
    .ZN(_0543_));
 XNOR2_X1 _4740_ (.A(_0488_),
    .B(_0543_),
    .ZN(_0544_));
 XOR2_X1 _4741_ (.A(_0487_),
    .B(_0544_),
    .Z(_0545_));
 XNOR2_X1 _4742_ (.A(_0486_),
    .B(_0545_),
    .ZN(_0546_));
 XNOR2_X1 _4743_ (.A(_0484_),
    .B(_0546_),
    .ZN(_0547_));
 XNOR2_X1 _4744_ (.A(_0480_),
    .B(_0547_),
    .ZN(_0548_));
 XNOR2_X1 _4745_ (.A(_0476_),
    .B(_0548_),
    .ZN(_0549_));
 XNOR2_X1 _4746_ (.A(_0474_),
    .B(_0549_),
    .ZN(_0550_));
 XOR2_X1 _4747_ (.A(_0462_),
    .B(_0550_),
    .Z(_0551_));
 XNOR2_X1 _4748_ (.A(_0460_),
    .B(_0551_),
    .ZN(_0552_));
 XOR2_X1 _4749_ (.A(_0444_),
    .B(_0552_),
    .Z(_0553_));
 XNOR2_X1 _4750_ (.A(_0442_),
    .B(_0553_),
    .ZN(_0554_));
 XOR2_X1 _4751_ (.A(_0439_),
    .B(_0554_),
    .Z(_0555_));
 XNOR2_X1 _4752_ (.A(_0437_),
    .B(_0555_),
    .ZN(_0556_));
 XNOR2_X1 _4753_ (.A(_0434_),
    .B(_0556_),
    .ZN(_0557_));
 XOR2_X1 _4754_ (.A(_0433_),
    .B(_0557_),
    .Z(_0558_));
 XNOR2_X1 _4755_ (.A(_0431_),
    .B(_0558_),
    .ZN(_0559_));
 XOR2_X1 _4756_ (.A(_0430_),
    .B(_0559_),
    .Z(_0560_));
 XNOR2_X1 _4757_ (.A(_0428_),
    .B(_0560_),
    .ZN(_0561_));
 NOR2_X1 _4758_ (.A1(_0426_),
    .A2(_0561_),
    .ZN(_0562_));
 XOR2_X1 _4759_ (.A(_0426_),
    .B(_0561_),
    .Z(_0563_));
 NOR2_X1 _4760_ (.A1(_0012_),
    .A2(_0423_),
    .ZN(_0564_));
 AOI21_X1 _4761_ (.A(_0562_),
    .B1(_0563_),
    .B2(_0564_),
    .ZN(_0565_));
 NOR2_X1 _4762_ (.A1(_0022_),
    .A2(_0427_),
    .ZN(_0566_));
 NOR2_X1 _4763_ (.A1(_0430_),
    .A2(_0559_),
    .ZN(_0567_));
 AOI21_X1 _4764_ (.A(_0567_),
    .B1(_0560_),
    .B2(_0428_),
    .ZN(_0568_));
 NAND2_X1 _4765_ (.A1(\fir.p5[8] ),
    .A2(\fir.p5[6] ),
    .ZN(_0569_));
 XOR2_X1 _4766_ (.A(_0027_),
    .B(_0569_),
    .Z(_0570_));
 NOR2_X1 _4767_ (.A1(_0433_),
    .A2(_0557_),
    .ZN(_0571_));
 AOI21_X1 _4768_ (.A(_0571_),
    .B1(_0558_),
    .B2(_0431_),
    .ZN(_0572_));
 XNOR2_X1 _4769_ (.A(\fir.p5[9] ),
    .B(\fir.p5[7] ),
    .ZN(_0573_));
 NOR2_X1 _4770_ (.A1(_0434_),
    .A2(_0556_),
    .ZN(_0574_));
 INV_X1 _4771_ (.A(\fir.p5[11] ),
    .ZN(_0575_));
 NOR2_X1 _4772_ (.A1(_0439_),
    .A2(_0554_),
    .ZN(_0576_));
 AOI21_X1 _4773_ (.A(_0576_),
    .B1(_0555_),
    .B2(_0437_),
    .ZN(_0577_));
 NOR2_X1 _4774_ (.A1(_0444_),
    .A2(_0552_),
    .ZN(_0578_));
 AOI21_X1 _4775_ (.A(_0578_),
    .B1(_0553_),
    .B2(_0442_),
    .ZN(_0579_));
 INV_X1 _4776_ (.A(_0457_),
    .ZN(_0580_));
 AOI21_X1 _4777_ (.A(_0580_),
    .B1(_0458_),
    .B2(_0446_),
    .ZN(_0581_));
 NAND2_X1 _4778_ (.A1(_0460_),
    .A2(_0551_),
    .ZN(_0582_));
 OAI21_X1 _4779_ (.A(_0582_),
    .B1(_0550_),
    .B2(_0462_),
    .ZN(_0583_));
 INV_X1 _4780_ (.A(_0453_),
    .ZN(_0584_));
 NOR2_X1 _4781_ (.A1(_0449_),
    .A2(_0584_),
    .ZN(_0585_));
 NOR2_X1 _4782_ (.A1(_3587_),
    .A2(_0451_),
    .ZN(_0586_));
 NOR2_X1 _4783_ (.A1(_3599_),
    .A2(_0452_),
    .ZN(_0587_));
 NOR2_X1 _4784_ (.A1(_0586_),
    .A2(_0587_),
    .ZN(_0588_));
 AND2_X1 _4785_ (.A1(\fir.p3[9] ),
    .A2(\fir.p3[8] ),
    .ZN(_0589_));
 AOI21_X1 _4786_ (.A(_0589_),
    .B1(_0466_),
    .B2(\fir.p3[7] ),
    .ZN(_0590_));
 XNOR2_X1 _4787_ (.A(_0254_),
    .B(_0590_),
    .ZN(_0591_));
 XOR2_X1 _4788_ (.A(_0267_),
    .B(_0591_),
    .Z(_0592_));
 XNOR2_X1 _4789_ (.A(_0588_),
    .B(_0592_),
    .ZN(_0593_));
 NOR2_X1 _4790_ (.A1(_0464_),
    .A2(_0472_),
    .ZN(_0594_));
 NOR2_X1 _4791_ (.A1(_0468_),
    .A2(_0471_),
    .ZN(_0595_));
 OAI21_X1 _4792_ (.A(_0593_),
    .B1(_0594_),
    .B2(_0595_),
    .ZN(_0596_));
 OR3_X1 _4793_ (.A1(_0595_),
    .A2(_0594_),
    .A3(_0593_),
    .ZN(_0597_));
 AND2_X1 _4794_ (.A1(_0596_),
    .A2(_0597_),
    .ZN(_0598_));
 XNOR2_X1 _4795_ (.A(_0585_),
    .B(_0598_),
    .ZN(_0599_));
 NAND2_X1 _4796_ (.A1(_0476_),
    .A2(_0548_),
    .ZN(_0600_));
 OAI21_X1 _4797_ (.A(_0600_),
    .B1(_0549_),
    .B2(_0474_),
    .ZN(_0601_));
 OR2_X1 _4798_ (.A1(_0465_),
    .A2(_0467_),
    .ZN(_0602_));
 XOR2_X1 _4799_ (.A(\fir.p3[9] ),
    .B(\fir.p3[10] ),
    .Z(_0603_));
 XNOR2_X1 _4800_ (.A(\fir.p3[8] ),
    .B(_0603_),
    .ZN(_0604_));
 XNOR2_X1 _4801_ (.A(_0465_),
    .B(_0604_),
    .ZN(_0605_));
 NOR2_X1 _4802_ (.A1(_3574_),
    .A2(_0478_),
    .ZN(_0606_));
 NOR2_X1 _4803_ (.A1(_3579_),
    .A2(_0479_),
    .ZN(_0607_));
 NOR2_X1 _4804_ (.A1(_0606_),
    .A2(_0607_),
    .ZN(_0608_));
 XNOR2_X1 _4805_ (.A(_0605_),
    .B(_0608_),
    .ZN(_0609_));
 XNOR2_X1 _4806_ (.A(_0602_),
    .B(_0609_),
    .ZN(_0610_));
 NAND2_X1 _4807_ (.A1(_0484_),
    .A2(_0546_),
    .ZN(_0611_));
 INV_X1 _4808_ (.A(_0480_),
    .ZN(_0612_));
 OAI21_X1 _4809_ (.A(_0611_),
    .B1(_0547_),
    .B2(_0612_),
    .ZN(_0613_));
 AND2_X1 _4810_ (.A1(\fir.p4[9] ),
    .A2(\fir.p4[8] ),
    .ZN(_0614_));
 AOI21_X1 _4811_ (.A(_0614_),
    .B1(_0485_),
    .B2(\fir.p4[7] ),
    .ZN(_0615_));
 XNOR2_X1 _4812_ (.A(_0242_),
    .B(_0615_),
    .ZN(_0616_));
 XOR2_X1 _4813_ (.A(_0246_),
    .B(_0616_),
    .Z(_0617_));
 INV_X1 _4814_ (.A(_0486_),
    .ZN(_0618_));
 NAND2_X1 _4815_ (.A1(_0618_),
    .A2(_0545_),
    .ZN(_0619_));
 OAI21_X1 _4816_ (.A(_0619_),
    .B1(_0544_),
    .B2(_0487_),
    .ZN(_0620_));
 OR2_X1 _4817_ (.A1(\fir.p4[9] ),
    .A2(\fir.p4[10] ),
    .ZN(_0621_));
 NAND2_X1 _4818_ (.A1(\fir.p4[9] ),
    .A2(\fir.p4[10] ),
    .ZN(_0622_));
 NAND2_X1 _4819_ (.A1(_0621_),
    .A2(_0622_),
    .ZN(_0623_));
 XNOR2_X1 _4820_ (.A(_3517_),
    .B(_0623_),
    .ZN(_0624_));
 NOR2_X1 _4821_ (.A1(_0026_),
    .A2(_0543_),
    .ZN(_0625_));
 NOR2_X1 _4822_ (.A1(_0494_),
    .A2(_0541_),
    .ZN(_0626_));
 AOI21_X1 _4823_ (.A(_0626_),
    .B1(_0542_),
    .B2(_0492_),
    .ZN(_0627_));
 NOR2_X1 _4824_ (.A1(_0498_),
    .A2(_0539_),
    .ZN(_0628_));
 AOI21_X1 _4825_ (.A(_0628_),
    .B1(_0540_),
    .B2(_0495_),
    .ZN(_0629_));
 NOR2_X1 _4826_ (.A1(_0019_),
    .A2(_0499_),
    .ZN(_0630_));
 NOR2_X1 _4827_ (.A1(_0503_),
    .A2(_0537_),
    .ZN(_0631_));
 AOI21_X1 _4828_ (.A(_0631_),
    .B1(_0538_),
    .B2(_0500_),
    .ZN(_0632_));
 NAND2_X1 _4829_ (.A1(\fir.p2[6] ),
    .A2(\fir.p2[10] ),
    .ZN(_0633_));
 XOR2_X1 _4830_ (.A(_0025_),
    .B(_0633_),
    .Z(_0634_));
 NOR2_X1 _4831_ (.A1(_0505_),
    .A2(_0535_),
    .ZN(_0635_));
 AOI21_X1 _4832_ (.A(_0635_),
    .B1(_0536_),
    .B2(_0504_),
    .ZN(_0636_));
 XOR2_X1 _4833_ (.A(\fir.p2[7] ),
    .B(\fir.p2[11] ),
    .Z(_0637_));
 NOR2_X1 _4834_ (.A1(_0024_),
    .A2(_0534_),
    .ZN(_0638_));
 NOR2_X1 _4835_ (.A1(_0510_),
    .A2(_0531_),
    .ZN(_0639_));
 NOR2_X1 _4836_ (.A1(_0513_),
    .A2(_0529_),
    .ZN(_0640_));
 AOI21_X1 _4837_ (.A(_0640_),
    .B1(_0530_),
    .B2(_0511_),
    .ZN(_0641_));
 NOR3_X1 _4838_ (.A1(\fir.p1[10] ),
    .A2(_0017_),
    .A3(_3663_),
    .ZN(_0642_));
 NOR2_X1 _4839_ (.A1(_0515_),
    .A2(_0527_),
    .ZN(_0643_));
 AOI21_X1 _4840_ (.A(_0643_),
    .B1(_0528_),
    .B2(_0514_),
    .ZN(_0644_));
 NOR2_X1 _4841_ (.A1(\fir.p1[11] ),
    .A2(_0374_),
    .ZN(_0645_));
 XNOR2_X1 _4842_ (.A(_0023_),
    .B(_0645_),
    .ZN(_0646_));
 NAND2_X1 _4843_ (.A1(\fir.p1[11] ),
    .A2(\fir.p1[10] ),
    .ZN(_0647_));
 NAND2_X1 _4844_ (.A1(\fir.p0[9] ),
    .A2(\fir.p0[11] ),
    .ZN(_0648_));
 XOR2_X1 _4845_ (.A(\fir.p0[11] ),
    .B(\fir.p0[10] ),
    .Z(_0649_));
 XNOR2_X1 _4846_ (.A(_0648_),
    .B(_0649_),
    .ZN(_0650_));
 XNOR2_X1 _4847_ (.A(\fir.p0[8] ),
    .B(_0650_),
    .ZN(_0651_));
 NAND2_X1 _4848_ (.A1(\fir.p0[7] ),
    .A2(_0520_),
    .ZN(_0652_));
 NAND3_X1 _4849_ (.A1(\fir.p0[8] ),
    .A2(\fir.p0[10] ),
    .A3(_0519_),
    .ZN(_0653_));
 AOI21_X1 _4850_ (.A(_0651_),
    .B1(_0652_),
    .B2(_0653_),
    .ZN(_0654_));
 AND3_X1 _4851_ (.A1(_0653_),
    .A2(_0652_),
    .A3(_0651_),
    .ZN(_0655_));
 OR2_X1 _4852_ (.A1(_0654_),
    .A2(_0655_),
    .ZN(_0656_));
 XOR2_X1 _4853_ (.A(_0647_),
    .B(_0656_),
    .Z(_0657_));
 NOR2_X1 _4854_ (.A1(_0517_),
    .A2(_0526_),
    .ZN(_0658_));
 OAI21_X1 _4855_ (.A(_0657_),
    .B1(_0658_),
    .B2(_0524_),
    .ZN(_0659_));
 OR3_X1 _4856_ (.A1(_0524_),
    .A2(_0658_),
    .A3(_0657_),
    .ZN(_0660_));
 AND2_X1 _4857_ (.A1(_0659_),
    .A2(_0660_),
    .ZN(_0661_));
 XNOR2_X1 _4858_ (.A(_0646_),
    .B(_0661_),
    .ZN(_0662_));
 XOR2_X1 _4859_ (.A(_0644_),
    .B(_0662_),
    .Z(_0663_));
 XNOR2_X1 _4860_ (.A(_0642_),
    .B(_0663_),
    .ZN(_0664_));
 XOR2_X1 _4861_ (.A(_0641_),
    .B(_0664_),
    .Z(_0665_));
 XNOR2_X1 _4862_ (.A(_0639_),
    .B(_0665_),
    .ZN(_0666_));
 NAND2_X1 _4863_ (.A1(_0508_),
    .A2(_0532_),
    .ZN(_0667_));
 OAI21_X1 _4864_ (.A(_0667_),
    .B1(_0533_),
    .B2(_0506_),
    .ZN(_0668_));
 NOR2_X1 _4865_ (.A1(_0393_),
    .A2(_0533_),
    .ZN(_0669_));
 NOR4_X1 _4866_ (.A1(_3557_),
    .A2(_0222_),
    .A3(_0393_),
    .A4(_0533_),
    .ZN(_0670_));
 AOI221_X1 _4867_ (.A(_0668_),
    .B1(_0669_),
    .B2(_0361_),
    .C1(_0670_),
    .C2(_3529_),
    .ZN(_0671_));
 XOR2_X1 _4868_ (.A(_0666_),
    .B(_0671_),
    .Z(_0672_));
 XNOR2_X1 _4869_ (.A(\fir.p2[9] ),
    .B(_0672_),
    .ZN(_0673_));
 XNOR2_X1 _4870_ (.A(_0638_),
    .B(_0673_),
    .ZN(_0674_));
 XNOR2_X1 _4871_ (.A(_0637_),
    .B(_0674_),
    .ZN(_0675_));
 XOR2_X1 _4872_ (.A(_0636_),
    .B(_0675_),
    .Z(_0676_));
 XNOR2_X1 _4873_ (.A(_0634_),
    .B(_0676_),
    .ZN(_0677_));
 XOR2_X1 _4874_ (.A(_0632_),
    .B(_0677_),
    .Z(_0678_));
 XNOR2_X1 _4875_ (.A(_0630_),
    .B(_0678_),
    .ZN(_0679_));
 XOR2_X1 _4876_ (.A(_0629_),
    .B(_0679_),
    .Z(_0680_));
 XOR2_X1 _4877_ (.A(_0627_),
    .B(_0680_),
    .Z(_0681_));
 XNOR2_X1 _4878_ (.A(\fir.p4[11] ),
    .B(_0681_),
    .ZN(_0682_));
 XNOR2_X1 _4879_ (.A(_0625_),
    .B(_0682_),
    .ZN(_0683_));
 XOR2_X1 _4880_ (.A(_0624_),
    .B(_0683_),
    .Z(_0684_));
 XNOR2_X1 _4881_ (.A(_0620_),
    .B(_0684_),
    .ZN(_0685_));
 XNOR2_X1 _4882_ (.A(_0617_),
    .B(_0685_),
    .ZN(_0686_));
 XOR2_X1 _4883_ (.A(_0613_),
    .B(_0686_),
    .Z(_0687_));
 XNOR2_X1 _4884_ (.A(_0610_),
    .B(_0687_),
    .ZN(_0688_));
 XNOR2_X1 _4885_ (.A(_0601_),
    .B(_0688_),
    .ZN(_0689_));
 XOR2_X1 _4886_ (.A(_0599_),
    .B(_0689_),
    .Z(_0690_));
 XNOR2_X1 _4887_ (.A(_0583_),
    .B(_0690_),
    .ZN(_0691_));
 XOR2_X1 _4888_ (.A(_0581_),
    .B(_0691_),
    .Z(_0692_));
 XNOR2_X1 _4889_ (.A(_0579_),
    .B(_0692_),
    .ZN(_0693_));
 XNOR2_X1 _4890_ (.A(_0577_),
    .B(_0693_),
    .ZN(_0694_));
 XNOR2_X1 _4891_ (.A(_0575_),
    .B(_0694_),
    .ZN(_0695_));
 XNOR2_X1 _4892_ (.A(_0574_),
    .B(_0695_),
    .ZN(_0696_));
 XNOR2_X1 _4893_ (.A(_0573_),
    .B(_0696_),
    .ZN(_0697_));
 XOR2_X1 _4894_ (.A(_0572_),
    .B(_0697_),
    .Z(_0698_));
 XNOR2_X1 _4895_ (.A(_0570_),
    .B(_0698_),
    .ZN(_0699_));
 XOR2_X1 _4896_ (.A(_0568_),
    .B(_0699_),
    .Z(_0700_));
 XNOR2_X1 _4897_ (.A(_0566_),
    .B(_0700_),
    .ZN(_0701_));
 OR2_X1 _4898_ (.A1(_0565_),
    .A2(_0701_),
    .ZN(_0702_));
 XNOR2_X1 _4899_ (.A(_0292_),
    .B(_0293_),
    .ZN(_0703_));
 XNOR2_X1 _4900_ (.A(\fir.p5[5] ),
    .B(\fir.p5[3] ),
    .ZN(_0704_));
 INV_X1 _4901_ (.A(net185),
    .ZN(_0705_));
 XNOR2_X1 _4902_ (.A(_3503_),
    .B(_3504_),
    .ZN(_0706_));
 NOR2_X1 _4903_ (.A1(_0705_),
    .A2(_0706_),
    .ZN(_0707_));
 XNOR2_X1 _4904_ (.A(\fir.p5[7] ),
    .B(_3619_),
    .ZN(_0708_));
 XOR2_X1 _4905_ (.A(_0707_),
    .B(_0708_),
    .Z(_0709_));
 OR2_X1 _4906_ (.A1(_0704_),
    .A2(_0709_),
    .ZN(_0710_));
 OR3_X1 _4907_ (.A1(_0705_),
    .A2(_0706_),
    .A3(_0708_),
    .ZN(_0711_));
 AOI21_X1 _4908_ (.A(_0703_),
    .B1(_0710_),
    .B2(_0711_),
    .ZN(_0712_));
 INV_X1 _4909_ (.A(_0712_),
    .ZN(_0713_));
 NAND2_X1 _4910_ (.A1(\fir.p5[5] ),
    .A2(\fir.p5[3] ),
    .ZN(_0714_));
 XOR2_X1 _4911_ (.A(_0013_),
    .B(_0714_),
    .Z(_0715_));
 INV_X1 _4912_ (.A(_0715_),
    .ZN(_0716_));
 NAND2_X1 _4913_ (.A1(_0711_),
    .A2(_0710_),
    .ZN(_0717_));
 XOR2_X1 _4914_ (.A(_0717_),
    .B(_0703_),
    .Z(_0718_));
 OAI21_X1 _4915_ (.A(_0713_),
    .B1(_0716_),
    .B2(_0718_),
    .ZN(_0719_));
 XOR2_X1 _4916_ (.A(_0424_),
    .B(_0425_),
    .Z(_0720_));
 NAND2_X1 _4917_ (.A1(_0719_),
    .A2(_0720_),
    .ZN(_0721_));
 XNOR2_X1 _4918_ (.A(_0719_),
    .B(_0720_),
    .ZN(_0722_));
 OR2_X1 _4919_ (.A1(_0013_),
    .A2(_0714_),
    .ZN(_0723_));
 OAI21_X1 _4920_ (.A(_0721_),
    .B1(_0722_),
    .B2(_0723_),
    .ZN(_0724_));
 XOR2_X1 _4921_ (.A(_0564_),
    .B(_0563_),
    .Z(_0725_));
 AND2_X1 _4922_ (.A1(_0724_),
    .A2(_0725_),
    .ZN(_0726_));
 NAND2_X1 _4923_ (.A1(\fir.p5[4] ),
    .A2(\fir.p5[2] ),
    .ZN(_0727_));
 NOR2_X1 _4924_ (.A1(_0014_),
    .A2(_0727_),
    .ZN(_0728_));
 AND3_X1 _4925_ (.A1(_3469_),
    .A2(_3479_),
    .A3(_3501_),
    .ZN(_0729_));
 NOR2_X1 _4926_ (.A1(_3502_),
    .A2(_0729_),
    .ZN(_0730_));
 NAND2_X1 _4927_ (.A1(\fir.p5[5] ),
    .A2(_0730_),
    .ZN(_0731_));
 XNOR2_X1 _4928_ (.A(_0705_),
    .B(_0706_),
    .ZN(_0732_));
 XOR2_X1 _4929_ (.A(_0731_),
    .B(_0732_),
    .Z(_0733_));
 XOR2_X1 _4930_ (.A(\fir.p5[4] ),
    .B(\fir.p5[2] ),
    .Z(_0734_));
 NAND2_X1 _4931_ (.A1(_0733_),
    .A2(_0734_),
    .ZN(_0735_));
 OAI21_X1 _4932_ (.A(_0735_),
    .B1(_0732_),
    .B2(_0731_),
    .ZN(_0736_));
 XOR2_X1 _4933_ (.A(_0704_),
    .B(_0709_),
    .Z(_0737_));
 NAND2_X1 _4934_ (.A1(_0736_),
    .A2(_0737_),
    .ZN(_0738_));
 XNOR2_X1 _4935_ (.A(_0736_),
    .B(_0737_),
    .ZN(_0739_));
 XOR2_X1 _4936_ (.A(_0014_),
    .B(_0727_),
    .Z(_0740_));
 INV_X1 _4937_ (.A(_0740_),
    .ZN(_0741_));
 OAI21_X1 _4938_ (.A(_0738_),
    .B1(_0739_),
    .B2(_0741_),
    .ZN(_0742_));
 XNOR2_X1 _4939_ (.A(_0716_),
    .B(_0718_),
    .ZN(_0743_));
 XNOR2_X1 _4940_ (.A(_0742_),
    .B(_0743_),
    .ZN(_0744_));
 NAND2_X1 _4941_ (.A1(_0728_),
    .A2(_0744_),
    .ZN(_0745_));
 INV_X1 _4942_ (.A(_0742_),
    .ZN(_0746_));
 OAI21_X1 _4943_ (.A(_0745_),
    .B1(_0743_),
    .B2(_0746_),
    .ZN(_0747_));
 XOR2_X1 _4944_ (.A(_0723_),
    .B(_0722_),
    .Z(_0748_));
 NAND2_X1 _4945_ (.A1(_0747_),
    .A2(_0748_),
    .ZN(_0749_));
 NOR2_X1 _4946_ (.A1(_0747_),
    .A2(_0748_),
    .ZN(_0750_));
 XNOR2_X1 _4947_ (.A(_3480_),
    .B(_3500_),
    .ZN(_0751_));
 NAND2_X1 _4948_ (.A1(\fir.p5[4] ),
    .A2(_0751_),
    .ZN(_0752_));
 XNOR2_X1 _4949_ (.A(\fir.p5[5] ),
    .B(_0730_),
    .ZN(_0753_));
 NOR2_X1 _4950_ (.A1(_0752_),
    .A2(_0753_),
    .ZN(_0754_));
 XOR2_X1 _4951_ (.A(\fir.p5[3] ),
    .B(\fir.p5[1] ),
    .Z(_0755_));
 XOR2_X1 _4952_ (.A(_0752_),
    .B(_0753_),
    .Z(_0756_));
 AOI21_X1 _4953_ (.A(_0754_),
    .B1(_0755_),
    .B2(_0756_),
    .ZN(_0757_));
 XNOR2_X1 _4954_ (.A(_0733_),
    .B(_0734_),
    .ZN(_0758_));
 NOR2_X1 _4955_ (.A1(_0757_),
    .A2(_0758_),
    .ZN(_0759_));
 NAND2_X1 _4956_ (.A1(\fir.p5[3] ),
    .A2(\fir.p5[1] ),
    .ZN(_0760_));
 XOR2_X1 _4957_ (.A(_0015_),
    .B(_0760_),
    .Z(_0761_));
 XOR2_X1 _4958_ (.A(_0757_),
    .B(_0758_),
    .Z(_0762_));
 AOI21_X1 _4959_ (.A(_0759_),
    .B1(_0761_),
    .B2(_0762_),
    .ZN(_0763_));
 XNOR2_X1 _4960_ (.A(_0739_),
    .B(_0740_),
    .ZN(_0764_));
 INV_X1 _4961_ (.A(_0764_),
    .ZN(_0765_));
 NOR2_X1 _4962_ (.A1(_0763_),
    .A2(_0765_),
    .ZN(_0766_));
 XNOR2_X1 _4963_ (.A(_0763_),
    .B(_0764_),
    .ZN(_0767_));
 NOR2_X1 _4964_ (.A1(_0015_),
    .A2(_0760_),
    .ZN(_0768_));
 AOI21_X1 _4965_ (.A(_0766_),
    .B1(_0767_),
    .B2(_0768_),
    .ZN(_0769_));
 XNOR2_X1 _4966_ (.A(_0728_),
    .B(_0744_),
    .ZN(_0770_));
 NOR2_X1 _4967_ (.A1(_0769_),
    .A2(_0770_),
    .ZN(_0771_));
 XOR2_X1 _4968_ (.A(_0755_),
    .B(_0756_),
    .Z(_0772_));
 XOR2_X1 _4969_ (.A(\fir.p5[2] ),
    .B(\fir.p5[0] ),
    .Z(_0773_));
 XNOR2_X1 _4970_ (.A(\fir.p5[4] ),
    .B(_0751_),
    .ZN(_0774_));
 XOR2_X1 _4971_ (.A(_3497_),
    .B(_3499_),
    .Z(_0775_));
 NAND2_X1 _4972_ (.A1(\fir.p5[3] ),
    .A2(_0775_),
    .ZN(_0776_));
 XOR2_X1 _4973_ (.A(_0774_),
    .B(_0776_),
    .Z(_0777_));
 AND2_X1 _4974_ (.A1(_0773_),
    .A2(_0777_),
    .ZN(_0778_));
 NOR2_X1 _4975_ (.A1(_0774_),
    .A2(_0776_),
    .ZN(_0779_));
 OAI21_X1 _4976_ (.A(_0772_),
    .B1(_0778_),
    .B2(_0779_),
    .ZN(_0780_));
 NOR2_X1 _4977_ (.A1(_0779_),
    .A2(_0778_),
    .ZN(_0781_));
 XNOR2_X1 _4978_ (.A(_0781_),
    .B(_0772_),
    .ZN(_0782_));
 NAND3_X1 _4979_ (.A1(\fir.p5[2] ),
    .A2(\fir.p5[0] ),
    .A3(_0782_),
    .ZN(_0783_));
 AND2_X1 _4980_ (.A1(_0780_),
    .A2(_0783_),
    .ZN(_0784_));
 XNOR2_X1 _4981_ (.A(_0761_),
    .B(_0762_),
    .ZN(_0785_));
 NOR2_X1 _4982_ (.A1(_0784_),
    .A2(_0785_),
    .ZN(_0786_));
 XOR2_X1 _4983_ (.A(_0768_),
    .B(_0767_),
    .Z(_0787_));
 NAND2_X1 _4984_ (.A1(_0786_),
    .A2(_0787_),
    .ZN(_0788_));
 NOR2_X1 _4985_ (.A1(_0786_),
    .A2(_0787_),
    .ZN(_0789_));
 NAND2_X1 _4986_ (.A1(\fir.p5[2] ),
    .A2(\fir.p5[0] ),
    .ZN(_0790_));
 XNOR2_X1 _4987_ (.A(_0790_),
    .B(_0782_),
    .ZN(_0791_));
 XNOR2_X1 _4988_ (.A(\fir.p5[3] ),
    .B(_0775_),
    .ZN(_0792_));
 NOR2_X1 _4989_ (.A1(_3487_),
    .A2(_3496_),
    .ZN(_0793_));
 XNOR2_X1 _4990_ (.A(_3488_),
    .B(_0793_),
    .ZN(_0794_));
 NAND2_X1 _4991_ (.A1(\fir.p5[2] ),
    .A2(_0794_),
    .ZN(_0795_));
 XOR2_X1 _4992_ (.A(_0792_),
    .B(_0795_),
    .Z(_0796_));
 XNOR2_X1 _4993_ (.A(\fir.p5[1] ),
    .B(_0796_),
    .ZN(_0797_));
 XNOR2_X1 _4994_ (.A(\fir.p5[2] ),
    .B(_0794_),
    .ZN(_0798_));
 XOR2_X1 _4995_ (.A(_3494_),
    .B(_3495_),
    .Z(_0799_));
 NAND2_X1 _4996_ (.A1(\fir.p5[1] ),
    .A2(_0799_),
    .ZN(_0800_));
 XOR2_X1 _4997_ (.A(_0798_),
    .B(_0800_),
    .Z(_0801_));
 NAND2_X1 _4998_ (.A1(\fir.p5[0] ),
    .A2(_0801_),
    .ZN(_0802_));
 OR2_X1 _4999_ (.A1(_0798_),
    .A2(_0800_),
    .ZN(_0803_));
 AOI21_X1 _5000_ (.A(_0797_),
    .B1(_0802_),
    .B2(_0803_),
    .ZN(_0804_));
 NAND2_X1 _5001_ (.A1(\fir.p5[1] ),
    .A2(_0796_),
    .ZN(_0805_));
 OAI21_X1 _5002_ (.A(_0805_),
    .B1(_0795_),
    .B2(_0792_),
    .ZN(_0806_));
 XOR2_X1 _5003_ (.A(_0773_),
    .B(_0777_),
    .Z(_0807_));
 XOR2_X1 _5004_ (.A(_0806_),
    .B(_0807_),
    .Z(_0808_));
 AND2_X1 _5005_ (.A1(_0804_),
    .A2(_0808_),
    .ZN(_0809_));
 XOR2_X1 _5006_ (.A(_3492_),
    .B(_3493_),
    .Z(_0810_));
 NAND2_X1 _5007_ (.A1(\fir.p5[0] ),
    .A2(_0810_),
    .ZN(_0811_));
 XNOR2_X1 _5008_ (.A(\fir.p5[1] ),
    .B(_0799_),
    .ZN(_0812_));
 XNOR2_X1 _5009_ (.A(\fir.p5[0] ),
    .B(_0801_),
    .ZN(_0813_));
 NOR3_X1 _5010_ (.A1(_0811_),
    .A2(_0812_),
    .A3(_0813_),
    .ZN(_0814_));
 AND3_X1 _5011_ (.A1(_0803_),
    .A2(_0802_),
    .A3(_0797_),
    .ZN(_0815_));
 NOR2_X1 _5012_ (.A1(_0804_),
    .A2(_0815_),
    .ZN(_0816_));
 NAND2_X1 _5013_ (.A1(_0814_),
    .A2(_0816_),
    .ZN(_0817_));
 XNOR2_X1 _5014_ (.A(_0804_),
    .B(_0808_),
    .ZN(_0818_));
 OR2_X1 _5015_ (.A1(_0817_),
    .A2(_0818_),
    .ZN(_0819_));
 INV_X1 _5016_ (.A(_0819_),
    .ZN(_0820_));
 AND2_X1 _5017_ (.A1(_0806_),
    .A2(_0807_),
    .ZN(_0821_));
 NOR2_X1 _5018_ (.A1(_0821_),
    .A2(_0809_),
    .ZN(_0822_));
 XNOR2_X1 _5019_ (.A(_0791_),
    .B(_0822_),
    .ZN(_0823_));
 AOI22_X1 _5020_ (.A1(_0791_),
    .A2(_0809_),
    .B1(_0820_),
    .B2(_0823_),
    .ZN(_0824_));
 XOR2_X1 _5021_ (.A(_0784_),
    .B(_0785_),
    .Z(_0825_));
 AND2_X1 _5022_ (.A1(_0821_),
    .A2(_0791_),
    .ZN(_0826_));
 XNOR2_X1 _5023_ (.A(_0825_),
    .B(_0826_),
    .ZN(_0827_));
 NOR2_X1 _5024_ (.A1(_0824_),
    .A2(_0827_),
    .ZN(_0828_));
 AOI21_X1 _5025_ (.A(_0828_),
    .B1(_0826_),
    .B2(_0825_),
    .ZN(_0829_));
 OAI21_X1 _5026_ (.A(_0788_),
    .B1(_0789_),
    .B2(_0829_),
    .ZN(_0830_));
 XOR2_X1 _5027_ (.A(_0769_),
    .B(_0770_),
    .Z(_0831_));
 AOI21_X1 _5028_ (.A(_0771_),
    .B1(_0830_),
    .B2(_0831_),
    .ZN(_0832_));
 OAI21_X1 _5029_ (.A(_0749_),
    .B1(_0750_),
    .B2(_0832_),
    .ZN(_0833_));
 OR2_X1 _5030_ (.A1(_0724_),
    .A2(_0725_),
    .ZN(_0834_));
 AOI21_X1 _5031_ (.A(_0726_),
    .B1(_0833_),
    .B2(_0834_),
    .ZN(_0835_));
 AND2_X1 _5032_ (.A1(_0565_),
    .A2(_0701_),
    .ZN(_0836_));
 OAI21_X1 _5033_ (.A(_0702_),
    .B1(_0835_),
    .B2(_0836_),
    .ZN(_0837_));
 NOR2_X1 _5034_ (.A1(_0568_),
    .A2(_0699_),
    .ZN(_0838_));
 AOI21_X1 _5035_ (.A(_0838_),
    .B1(_0700_),
    .B2(_0566_),
    .ZN(_0839_));
 OR2_X1 _5036_ (.A1(_0027_),
    .A2(_0569_),
    .ZN(_0840_));
 NOR2_X1 _5037_ (.A1(_0572_),
    .A2(_0697_),
    .ZN(_0841_));
 AOI21_X1 _5038_ (.A(_0841_),
    .B1(_0698_),
    .B2(_0570_),
    .ZN(_0842_));
 NAND2_X1 _5039_ (.A1(\fir.p5[9] ),
    .A2(\fir.p5[7] ),
    .ZN(_0843_));
 XOR2_X1 _5040_ (.A(_0030_),
    .B(_0843_),
    .Z(_0844_));
 NAND2_X1 _5041_ (.A1(_0574_),
    .A2(_0695_),
    .ZN(_0845_));
 OAI21_X1 _5042_ (.A(_0845_),
    .B1(_0696_),
    .B2(_0573_),
    .ZN(_0846_));
 XNOR2_X1 _5043_ (.A(\fir.p5[8] ),
    .B(\fir.p5[10] ),
    .ZN(_0847_));
 INV_X1 _5044_ (.A(_0029_),
    .ZN(_0848_));
 AND2_X1 _5045_ (.A1(_0848_),
    .A2(_0694_),
    .ZN(_0849_));
 NAND2_X1 _5046_ (.A1(_0583_),
    .A2(_0690_),
    .ZN(_0850_));
 OAI21_X1 _5047_ (.A(_0850_),
    .B1(_0691_),
    .B2(_0581_),
    .ZN(_0851_));
 NAND2_X1 _5048_ (.A1(_0585_),
    .A2(_0598_),
    .ZN(_0852_));
 NAND2_X1 _5049_ (.A1(_0596_),
    .A2(_0852_),
    .ZN(_0853_));
 NAND2_X1 _5050_ (.A1(_0601_),
    .A2(_0688_),
    .ZN(_0854_));
 OAI21_X1 _5051_ (.A(_0854_),
    .B1(_0689_),
    .B2(_0599_),
    .ZN(_0855_));
 INV_X1 _5052_ (.A(_0592_),
    .ZN(_0856_));
 NOR2_X1 _5053_ (.A1(_0588_),
    .A2(_0856_),
    .ZN(_0857_));
 NAND2_X1 _5054_ (.A1(\fir.p3[9] ),
    .A2(\fir.p3[10] ),
    .ZN(_0858_));
 NAND2_X1 _5055_ (.A1(\fir.p3[8] ),
    .A2(_0603_),
    .ZN(_0859_));
 AOI21_X1 _5056_ (.A(_0328_),
    .B1(_0858_),
    .B2(_0859_),
    .ZN(_0860_));
 AND3_X1 _5057_ (.A1(_0328_),
    .A2(_0858_),
    .A3(_0859_),
    .ZN(_0861_));
 OR2_X1 _5058_ (.A1(_0860_),
    .A2(_0861_),
    .ZN(_0862_));
 XOR2_X1 _5059_ (.A(_0314_),
    .B(_0862_),
    .Z(_0863_));
 NOR2_X1 _5060_ (.A1(_0267_),
    .A2(_0591_),
    .ZN(_0864_));
 NOR2_X1 _5061_ (.A1(_0254_),
    .A2(_0590_),
    .ZN(_0865_));
 OAI21_X1 _5062_ (.A(_0863_),
    .B1(_0864_),
    .B2(_0865_),
    .ZN(_0866_));
 OR3_X1 _5063_ (.A1(_0865_),
    .A2(_0864_),
    .A3(_0863_),
    .ZN(_0867_));
 AND2_X1 _5064_ (.A1(_0866_),
    .A2(_0867_),
    .ZN(_0868_));
 NOR2_X1 _5065_ (.A1(_0602_),
    .A2(_0609_),
    .ZN(_0869_));
 NOR2_X1 _5066_ (.A1(_0605_),
    .A2(_0608_),
    .ZN(_0870_));
 OAI21_X1 _5067_ (.A(_0868_),
    .B1(_0869_),
    .B2(_0870_),
    .ZN(_0871_));
 OR3_X1 _5068_ (.A1(_0870_),
    .A2(_0869_),
    .A3(_0868_),
    .ZN(_0872_));
 AND2_X1 _5069_ (.A1(_0871_),
    .A2(_0872_),
    .ZN(_0873_));
 XNOR2_X1 _5070_ (.A(_0857_),
    .B(_0873_),
    .ZN(_0874_));
 NAND2_X1 _5071_ (.A1(_0613_),
    .A2(_0686_),
    .ZN(_0875_));
 NOR2_X1 _5072_ (.A1(_0613_),
    .A2(_0686_),
    .ZN(_0876_));
 OAI21_X1 _5073_ (.A(_0875_),
    .B1(_0876_),
    .B2(_0610_),
    .ZN(_0877_));
 OR2_X1 _5074_ (.A1(_0465_),
    .A2(_0604_),
    .ZN(_0878_));
 NOR2_X1 _5075_ (.A1(_0242_),
    .A2(_0615_),
    .ZN(_0879_));
 NOR2_X1 _5076_ (.A1(_0246_),
    .A2(_0616_),
    .ZN(_0880_));
 NOR2_X1 _5077_ (.A1(_0879_),
    .A2(_0880_),
    .ZN(_0881_));
 XNOR2_X1 _5078_ (.A(_0603_),
    .B(_0881_),
    .ZN(_0882_));
 XNOR2_X1 _5079_ (.A(_0878_),
    .B(_0882_),
    .ZN(_0883_));
 NAND2_X1 _5080_ (.A1(_0620_),
    .A2(_0684_),
    .ZN(_0884_));
 INV_X1 _5081_ (.A(_0617_),
    .ZN(_0885_));
 OAI21_X1 _5082_ (.A(_0884_),
    .B1(_0685_),
    .B2(_0885_),
    .ZN(_0886_));
 NAND3_X1 _5083_ (.A1(\fir.p4[8] ),
    .A2(_0621_),
    .A3(_0622_),
    .ZN(_0887_));
 AOI21_X1 _5084_ (.A(_0346_),
    .B1(_0622_),
    .B2(_0887_),
    .ZN(_0888_));
 AND3_X1 _5085_ (.A1(_0346_),
    .A2(_0622_),
    .A3(_0887_),
    .ZN(_0889_));
 OR2_X1 _5086_ (.A1(_0888_),
    .A2(_0889_),
    .ZN(_0890_));
 XOR2_X1 _5087_ (.A(_0339_),
    .B(_0890_),
    .Z(_0891_));
 INV_X1 _5088_ (.A(_0891_),
    .ZN(_0892_));
 NAND2_X1 _5089_ (.A1(_0625_),
    .A2(_0682_),
    .ZN(_0893_));
 OAI21_X1 _5090_ (.A(_0893_),
    .B1(_0683_),
    .B2(_0624_),
    .ZN(_0894_));
 OR2_X1 _5091_ (.A1(\fir.p4[11] ),
    .A2(\fir.p4[10] ),
    .ZN(_0895_));
 NAND2_X1 _5092_ (.A1(\fir.p4[11] ),
    .A2(\fir.p4[10] ),
    .ZN(_0896_));
 NAND2_X1 _5093_ (.A1(_0895_),
    .A2(_0896_),
    .ZN(_0897_));
 XOR2_X1 _5094_ (.A(\fir.p4[9] ),
    .B(_0897_),
    .Z(_0898_));
 NOR2_X1 _5095_ (.A1(_0026_),
    .A2(_0681_),
    .ZN(_0899_));
 NAND3_X1 _5096_ (.A1(_0491_),
    .A2(_0542_),
    .A3(_0680_),
    .ZN(_0900_));
 NOR2_X1 _5097_ (.A1(_0629_),
    .A2(_0679_),
    .ZN(_0901_));
 AOI21_X1 _5098_ (.A(_0901_),
    .B1(_0680_),
    .B2(_0626_),
    .ZN(_0902_));
 NOR2_X1 _5099_ (.A1(_0237_),
    .A2(_0402_),
    .ZN(_0903_));
 NAND3_X1 _5100_ (.A1(_0903_),
    .A2(_0542_),
    .A3(_0680_),
    .ZN(_0904_));
 OAI211_X1 _5101_ (.A(_0900_),
    .B(_0902_),
    .C1(_3636_),
    .C2(_0904_),
    .ZN(_0905_));
 NOR2_X1 _5102_ (.A1(_0632_),
    .A2(_0677_),
    .ZN(_0906_));
 AOI21_X1 _5103_ (.A(_0906_),
    .B1(_0678_),
    .B2(_0630_),
    .ZN(_0907_));
 NOR2_X1 _5104_ (.A1(_0025_),
    .A2(_0633_),
    .ZN(_0908_));
 NOR2_X1 _5105_ (.A1(_0636_),
    .A2(_0675_),
    .ZN(_0909_));
 AOI21_X1 _5106_ (.A(_0909_),
    .B1(_0676_),
    .B2(_0634_),
    .ZN(_0910_));
 NAND2_X1 _5107_ (.A1(\fir.p2[7] ),
    .A2(\fir.p2[11] ),
    .ZN(_0911_));
 XOR2_X1 _5108_ (.A(_0005_),
    .B(_0911_),
    .Z(_0912_));
 NOR3_X1 _5109_ (.A1(_0024_),
    .A2(_0534_),
    .A3(_0673_),
    .ZN(_0913_));
 AOI21_X1 _5110_ (.A(_0913_),
    .B1(_0674_),
    .B2(_0637_),
    .ZN(_0914_));
 XOR2_X1 _5111_ (.A(\fir.p2[8] ),
    .B(\fir.p2[11] ),
    .Z(_0915_));
 NAND2_X1 _5112_ (.A1(\fir.p2[9] ),
    .A2(_0672_),
    .ZN(_0916_));
 NOR2_X1 _5113_ (.A1(_0641_),
    .A2(_0664_),
    .ZN(_0917_));
 NOR3_X1 _5114_ (.A1(\fir.p1[11] ),
    .A2(_0023_),
    .A3(_0374_),
    .ZN(_0918_));
 NOR2_X1 _5115_ (.A1(_0647_),
    .A2(_0656_),
    .ZN(_0919_));
 NOR2_X1 _5116_ (.A1(_0654_),
    .A2(_0919_),
    .ZN(_0920_));
 INV_X1 _5117_ (.A(net265),
    .ZN(_0921_));
 NAND2_X1 _5118_ (.A1(\fir.p0[8] ),
    .A2(_0650_),
    .ZN(_0922_));
 OAI21_X1 _5119_ (.A(_0922_),
    .B1(_0648_),
    .B2(\fir.p0[10] ),
    .ZN(_0923_));
 NAND2_X1 _5120_ (.A1(\fir.p0[11] ),
    .A2(\fir.p0[10] ),
    .ZN(_0924_));
 XOR2_X1 _5121_ (.A(_0028_),
    .B(_0924_),
    .Z(_0925_));
 XNOR2_X1 _5122_ (.A(_0923_),
    .B(_0925_),
    .ZN(_0926_));
 XNOR2_X1 _5123_ (.A(_0921_),
    .B(_0926_),
    .ZN(_0927_));
 XOR2_X1 _5124_ (.A(_0920_),
    .B(_0927_),
    .Z(_0928_));
 XNOR2_X1 _5125_ (.A(\fir.p1[7] ),
    .B(_0928_),
    .ZN(_0929_));
 NAND2_X1 _5126_ (.A1(_0646_),
    .A2(_0661_),
    .ZN(_0930_));
 AOI21_X1 _5127_ (.A(_0929_),
    .B1(_0930_),
    .B2(_0659_),
    .ZN(_0931_));
 AND3_X1 _5128_ (.A1(_0659_),
    .A2(_0930_),
    .A3(_0929_),
    .ZN(_0932_));
 NOR2_X1 _5129_ (.A1(_0931_),
    .A2(_0932_),
    .ZN(_0933_));
 XNOR2_X1 _5130_ (.A(_0918_),
    .B(_0933_),
    .ZN(_0934_));
 NAND2_X1 _5131_ (.A1(_0642_),
    .A2(_0663_),
    .ZN(_0935_));
 OR2_X1 _5132_ (.A1(_0644_),
    .A2(_0662_),
    .ZN(_0936_));
 AOI21_X1 _5133_ (.A(_0934_),
    .B1(_0935_),
    .B2(_0936_),
    .ZN(_0937_));
 AND3_X1 _5134_ (.A1(_0936_),
    .A2(_0935_),
    .A3(_0934_),
    .ZN(_0938_));
 NOR2_X1 _5135_ (.A1(_0937_),
    .A2(_0938_),
    .ZN(_0939_));
 XNOR2_X1 _5136_ (.A(_0917_),
    .B(_0939_),
    .ZN(_0940_));
 NAND2_X1 _5137_ (.A1(_0639_),
    .A2(_0665_),
    .ZN(_0941_));
 OR2_X1 _5138_ (.A1(_0666_),
    .A2(_0671_),
    .ZN(_0942_));
 NAND2_X1 _5139_ (.A1(_0941_),
    .A2(_0942_),
    .ZN(_0943_));
 XNOR2_X1 _5140_ (.A(_0940_),
    .B(_0943_),
    .ZN(_0944_));
 XNOR2_X1 _5141_ (.A(\fir.p2[10] ),
    .B(_0944_),
    .ZN(_0945_));
 XOR2_X1 _5142_ (.A(_0916_),
    .B(_0945_),
    .Z(_0946_));
 XNOR2_X1 _5143_ (.A(_0915_),
    .B(_0946_),
    .ZN(_0947_));
 XOR2_X1 _5144_ (.A(_0914_),
    .B(_0947_),
    .Z(_0948_));
 XNOR2_X1 _5145_ (.A(_0912_),
    .B(_0948_),
    .ZN(_0949_));
 XOR2_X1 _5146_ (.A(_0910_),
    .B(_0949_),
    .Z(_0950_));
 XOR2_X1 _5147_ (.A(_0908_),
    .B(_0950_),
    .Z(_0951_));
 XNOR2_X1 _5148_ (.A(_0907_),
    .B(_0951_),
    .ZN(_0952_));
 XOR2_X1 _5149_ (.A(_0905_),
    .B(_0952_),
    .Z(_0953_));
 XNOR2_X1 _5150_ (.A(\fir.p4[11] ),
    .B(_0953_),
    .ZN(_0954_));
 XOR2_X1 _5151_ (.A(_0899_),
    .B(_0954_),
    .Z(_0955_));
 XOR2_X1 _5152_ (.A(_0898_),
    .B(_0955_),
    .Z(_0956_));
 XNOR2_X1 _5153_ (.A(_0894_),
    .B(_0956_),
    .ZN(_0957_));
 XNOR2_X1 _5154_ (.A(_0892_),
    .B(_0957_),
    .ZN(_0958_));
 XOR2_X1 _5155_ (.A(_0886_),
    .B(_0958_),
    .Z(_0959_));
 XNOR2_X1 _5156_ (.A(_0883_),
    .B(_0959_),
    .ZN(_0960_));
 XOR2_X1 _5157_ (.A(_0877_),
    .B(_0960_),
    .Z(_0961_));
 XNOR2_X1 _5158_ (.A(_0874_),
    .B(_0961_),
    .ZN(_0962_));
 XNOR2_X1 _5159_ (.A(_0855_),
    .B(_0962_),
    .ZN(_0963_));
 XNOR2_X1 _5160_ (.A(_0853_),
    .B(_0963_),
    .ZN(_0964_));
 XOR2_X1 _5161_ (.A(_0851_),
    .B(_0964_),
    .Z(_0965_));
 INV_X1 _5162_ (.A(_0579_),
    .ZN(_0966_));
 NAND2_X1 _5163_ (.A1(_0966_),
    .A2(_0692_),
    .ZN(_0967_));
 NOR2_X1 _5164_ (.A1(_0966_),
    .A2(_0692_),
    .ZN(_0968_));
 OAI21_X1 _5165_ (.A(_0967_),
    .B1(_0968_),
    .B2(_0577_),
    .ZN(_0969_));
 XNOR2_X1 _5166_ (.A(_0965_),
    .B(_0969_),
    .ZN(_0970_));
 XNOR2_X1 _5167_ (.A(\fir.p5[11] ),
    .B(_0970_),
    .ZN(_0971_));
 XOR2_X1 _5168_ (.A(_0849_),
    .B(_0971_),
    .Z(_0972_));
 XNOR2_X1 _5169_ (.A(_0847_),
    .B(_0972_),
    .ZN(_0973_));
 XOR2_X1 _5170_ (.A(_0846_),
    .B(_0973_),
    .Z(_0974_));
 XNOR2_X1 _5171_ (.A(_0844_),
    .B(_0974_),
    .ZN(_0975_));
 XOR2_X1 _5172_ (.A(_0842_),
    .B(_0975_),
    .Z(_0976_));
 XOR2_X1 _5173_ (.A(_0840_),
    .B(_0976_),
    .Z(_0977_));
 XOR2_X1 _5174_ (.A(_0839_),
    .B(_0977_),
    .Z(_0978_));
 XOR2_X1 _5175_ (.A(_0837_),
    .B(_0978_),
    .Z(_0979_));
 XOR2_X1 _5176_ (.A(_0565_),
    .B(_0701_),
    .Z(_0980_));
 XNOR2_X1 _5177_ (.A(_0835_),
    .B(_0980_),
    .ZN(_0981_));
 NAND2_X1 _5178_ (.A1(\fir.p7[11] ),
    .A2(_0981_),
    .ZN(_0982_));
 NOR2_X1 _5179_ (.A1(_0979_),
    .A2(_0982_),
    .ZN(_0983_));
 INV_X1 _5180_ (.A(\fir.p7[11] ),
    .ZN(_0984_));
 NOR2_X1 _5181_ (.A1(_0984_),
    .A2(_0981_),
    .ZN(_0985_));
 XNOR2_X1 _5182_ (.A(_0979_),
    .B(_0985_),
    .ZN(_0986_));
 INV_X1 _5183_ (.A(_0986_),
    .ZN(_0987_));
 XOR2_X1 _5184_ (.A(\fir.p7[11] ),
    .B(\fir.p7[9] ),
    .Z(_0988_));
 AOI21_X1 _5185_ (.A(_0983_),
    .B1(_0987_),
    .B2(_0988_),
    .ZN(_0989_));
 XOR2_X1 _5186_ (.A(\fir.p7[11] ),
    .B(\fir.p7[10] ),
    .Z(_0990_));
 INV_X1 _5187_ (.A(_0016_),
    .ZN(_0991_));
 AND2_X1 _5188_ (.A1(_0991_),
    .A2(_0979_),
    .ZN(_0992_));
 OR2_X1 _5189_ (.A1(_0842_),
    .A2(_0975_),
    .ZN(_0993_));
 AND2_X1 _5190_ (.A1(_0842_),
    .A2(_0975_),
    .ZN(_0994_));
 OAI21_X1 _5191_ (.A(_0993_),
    .B1(_0994_),
    .B2(_0840_),
    .ZN(_0995_));
 NOR2_X1 _5192_ (.A1(_0030_),
    .A2(_0843_),
    .ZN(_0996_));
 NAND2_X1 _5193_ (.A1(_0846_),
    .A2(_0973_),
    .ZN(_0997_));
 NOR2_X1 _5194_ (.A1(_0846_),
    .A2(_0973_),
    .ZN(_0998_));
 INV_X1 _5195_ (.A(_0844_),
    .ZN(_0999_));
 OAI21_X1 _5196_ (.A(_0997_),
    .B1(_0998_),
    .B2(_0999_),
    .ZN(_1000_));
 NAND2_X1 _5197_ (.A1(\fir.p5[8] ),
    .A2(\fir.p5[10] ),
    .ZN(_1001_));
 XOR2_X1 _5198_ (.A(_0033_),
    .B(_1001_),
    .Z(_1002_));
 NAND2_X1 _5199_ (.A1(_0849_),
    .A2(_0971_),
    .ZN(_1003_));
 NOR2_X1 _5200_ (.A1(_0849_),
    .A2(_0971_),
    .ZN(_1004_));
 OAI21_X1 _5201_ (.A(_1003_),
    .B1(_1004_),
    .B2(_0847_),
    .ZN(_1005_));
 XOR2_X1 _5202_ (.A(\fir.p5[9] ),
    .B(\fir.p5[11] ),
    .Z(_1006_));
 NOR2_X1 _5203_ (.A1(_0029_),
    .A2(_0970_),
    .ZN(_1007_));
 AOI21_X1 _5204_ (.A(_0963_),
    .B1(_0852_),
    .B2(_0596_),
    .ZN(_1008_));
 AOI21_X1 _5205_ (.A(_1008_),
    .B1(_0962_),
    .B2(_0855_),
    .ZN(_1009_));
 NAND2_X1 _5206_ (.A1(_0857_),
    .A2(_0873_),
    .ZN(_1010_));
 NAND2_X1 _5207_ (.A1(_0871_),
    .A2(_1010_),
    .ZN(_1011_));
 NAND2_X1 _5208_ (.A1(_0877_),
    .A2(_0960_),
    .ZN(_1012_));
 NOR2_X1 _5209_ (.A1(_0877_),
    .A2(_0960_),
    .ZN(_1013_));
 OAI21_X1 _5210_ (.A(_1012_),
    .B1(_1013_),
    .B2(_0874_),
    .ZN(_1014_));
 INV_X1 _5211_ (.A(_0860_),
    .ZN(_1015_));
 OAI21_X1 _5212_ (.A(_1015_),
    .B1(_0861_),
    .B2(_0314_),
    .ZN(_1016_));
 OAI21_X1 _5213_ (.A(\fir.p3[11] ),
    .B1(\fir.p3[10] ),
    .B2(\fir.p3[9] ),
    .ZN(_1017_));
 AND2_X1 _5214_ (.A1(_0858_),
    .A2(_1017_),
    .ZN(_1018_));
 XNOR2_X1 _5215_ (.A(_0467_),
    .B(_1018_),
    .ZN(_1019_));
 XOR2_X1 _5216_ (.A(_0451_),
    .B(_1019_),
    .Z(_1020_));
 XNOR2_X1 _5217_ (.A(_1016_),
    .B(_1020_),
    .ZN(_1021_));
 INV_X1 _5218_ (.A(_0881_),
    .ZN(_1022_));
 INV_X1 _5219_ (.A(_0878_),
    .ZN(_1023_));
 AOI22_X1 _5220_ (.A1(_0603_),
    .A2(_1022_),
    .B1(_0882_),
    .B2(_1023_),
    .ZN(_1024_));
 XNOR2_X1 _5221_ (.A(_1021_),
    .B(_1024_),
    .ZN(_1025_));
 XNOR2_X1 _5222_ (.A(_0866_),
    .B(_1025_),
    .ZN(_1026_));
 INV_X1 _5223_ (.A(_0958_),
    .ZN(_1027_));
 NAND2_X1 _5224_ (.A1(_0886_),
    .A2(_1027_),
    .ZN(_1028_));
 INV_X1 _5225_ (.A(_0883_),
    .ZN(_1029_));
 OAI21_X1 _5226_ (.A(_1028_),
    .B1(_0959_),
    .B2(_1029_),
    .ZN(_1030_));
 OR2_X1 _5227_ (.A1(_0465_),
    .A2(_0603_),
    .ZN(_1031_));
 XOR2_X1 _5228_ (.A(\fir.p3[11] ),
    .B(\fir.p3[10] ),
    .Z(_1032_));
 INV_X1 _5229_ (.A(_0888_),
    .ZN(_1033_));
 OAI21_X1 _5230_ (.A(_1033_),
    .B1(_0889_),
    .B2(_0339_),
    .ZN(_1034_));
 XNOR2_X1 _5231_ (.A(_1032_),
    .B(_1034_),
    .ZN(_1035_));
 XNOR2_X1 _5232_ (.A(_1031_),
    .B(_1035_),
    .ZN(_1036_));
 NAND2_X1 _5233_ (.A1(_0894_),
    .A2(_0956_),
    .ZN(_1037_));
 OAI21_X1 _5234_ (.A(_1037_),
    .B1(_0957_),
    .B2(_0892_),
    .ZN(_1038_));
 INV_X1 _5235_ (.A(_0896_),
    .ZN(_1039_));
 AOI21_X1 _5236_ (.A(_1039_),
    .B1(_0895_),
    .B2(\fir.p4[9] ),
    .ZN(_1040_));
 XNOR2_X1 _5237_ (.A(_0486_),
    .B(_1040_),
    .ZN(_1041_));
 XOR2_X1 _5238_ (.A(_0478_),
    .B(_1041_),
    .Z(_1042_));
 NOR3_X1 _5239_ (.A1(_0026_),
    .A2(_0681_),
    .A3(_0954_),
    .ZN(_1043_));
 NOR2_X1 _5240_ (.A1(_0898_),
    .A2(_0955_),
    .ZN(_1044_));
 NOR2_X1 _5241_ (.A1(_1043_),
    .A2(_1044_),
    .ZN(_1045_));
 INV_X1 _5242_ (.A(_0026_),
    .ZN(_1046_));
 NAND2_X1 _5243_ (.A1(_1046_),
    .A2(_0953_),
    .ZN(_1047_));
 NAND2_X1 _5244_ (.A1(_0908_),
    .A2(_0950_),
    .ZN(_1048_));
 OAI21_X1 _5245_ (.A(_1048_),
    .B1(_0949_),
    .B2(_0910_),
    .ZN(_1049_));
 NOR2_X1 _5246_ (.A1(_0005_),
    .A2(_0911_),
    .ZN(_1050_));
 NOR2_X1 _5247_ (.A1(_0914_),
    .A2(_0947_),
    .ZN(_1051_));
 AOI21_X1 _5248_ (.A(_1051_),
    .B1(_0948_),
    .B2(_0912_),
    .ZN(_1052_));
 NAND2_X1 _5249_ (.A1(\fir.p2[8] ),
    .A2(\fir.p2[11] ),
    .ZN(_1053_));
 XOR2_X1 _5250_ (.A(_0018_),
    .B(_1053_),
    .Z(_1054_));
 NAND2_X1 _5251_ (.A1(_0915_),
    .A2(_0946_),
    .ZN(_1055_));
 OAI21_X1 _5252_ (.A(_1055_),
    .B1(_0945_),
    .B2(_0916_),
    .ZN(_1056_));
 XOR2_X1 _5253_ (.A(\fir.p2[9] ),
    .B(\fir.p2[11] ),
    .Z(_1057_));
 AND2_X1 _5254_ (.A1(\fir.p2[10] ),
    .A2(_0944_),
    .ZN(_1058_));
 NOR2_X1 _5255_ (.A1(_0920_),
    .A2(_0927_),
    .ZN(_1059_));
 AOI21_X1 _5256_ (.A(_1059_),
    .B1(_0928_),
    .B2(\fir.p1[7] ),
    .ZN(_1060_));
 NOR2_X1 _5257_ (.A1(_0028_),
    .A2(_0924_),
    .ZN(_1061_));
 OAI21_X1 _5258_ (.A(\fir.p1[11] ),
    .B1(_0649_),
    .B2(_1061_),
    .ZN(_1062_));
 OR3_X1 _5259_ (.A1(\fir.p1[11] ),
    .A2(_0649_),
    .A3(_1061_),
    .ZN(_1063_));
 AND2_X1 _5260_ (.A1(_1062_),
    .A2(_1063_),
    .ZN(_1064_));
 NOR2_X1 _5261_ (.A1(_0921_),
    .A2(_0926_),
    .ZN(_1065_));
 AND2_X1 _5262_ (.A1(_0923_),
    .A2(_0925_),
    .ZN(_1066_));
 OAI21_X1 _5263_ (.A(_1064_),
    .B1(_1065_),
    .B2(_1066_),
    .ZN(_1067_));
 OR3_X1 _5264_ (.A1(_1066_),
    .A2(_1065_),
    .A3(_1064_),
    .ZN(_1068_));
 AND2_X1 _5265_ (.A1(_1067_),
    .A2(_1068_),
    .ZN(_1069_));
 XNOR2_X1 _5266_ (.A(\fir.p1[8] ),
    .B(_1069_),
    .ZN(_1070_));
 XOR2_X1 _5267_ (.A(_1060_),
    .B(_1070_),
    .Z(_1071_));
 AND2_X1 _5268_ (.A1(_0918_),
    .A2(_0933_),
    .ZN(_1072_));
 OAI21_X1 _5269_ (.A(_1071_),
    .B1(_1072_),
    .B2(_0931_),
    .ZN(_1073_));
 OR3_X1 _5270_ (.A1(_0931_),
    .A2(_1072_),
    .A3(_1071_),
    .ZN(_1074_));
 AND2_X1 _5271_ (.A1(_1073_),
    .A2(_1074_),
    .ZN(_1075_));
 XNOR2_X1 _5272_ (.A(_0937_),
    .B(_1075_),
    .ZN(_1076_));
 INV_X1 _5273_ (.A(_1076_),
    .ZN(_1077_));
 NAND2_X1 _5274_ (.A1(_0917_),
    .A2(_0939_),
    .ZN(_1078_));
 OAI21_X1 _5275_ (.A(_1078_),
    .B1(_0940_),
    .B2(_0941_),
    .ZN(_1079_));
 NOR2_X1 _5276_ (.A1(_0942_),
    .A2(_0940_),
    .ZN(_1080_));
 OAI21_X1 _5277_ (.A(_1077_),
    .B1(_1079_),
    .B2(_1080_),
    .ZN(_1081_));
 OR3_X1 _5278_ (.A1(_1080_),
    .A2(_1079_),
    .A3(_1077_),
    .ZN(_1082_));
 AND2_X1 _5279_ (.A1(_1081_),
    .A2(_1082_),
    .ZN(_1083_));
 XNOR2_X1 _5280_ (.A(\fir.p2[11] ),
    .B(_1083_),
    .ZN(_1084_));
 XNOR2_X1 _5281_ (.A(_1058_),
    .B(_1084_),
    .ZN(_1085_));
 XOR2_X1 _5282_ (.A(_1057_),
    .B(_1085_),
    .Z(_1086_));
 XOR2_X1 _5283_ (.A(_1056_),
    .B(_1086_),
    .Z(_1087_));
 XNOR2_X1 _5284_ (.A(_1054_),
    .B(_1087_),
    .ZN(_1088_));
 XOR2_X1 _5285_ (.A(_1052_),
    .B(_1088_),
    .Z(_1089_));
 XOR2_X1 _5286_ (.A(_1050_),
    .B(_1089_),
    .Z(_1090_));
 XNOR2_X1 _5287_ (.A(_1049_),
    .B(_1090_),
    .ZN(_1091_));
 INV_X1 _5288_ (.A(_0907_),
    .ZN(_1092_));
 AND2_X1 _5289_ (.A1(_1092_),
    .A2(_0951_),
    .ZN(_1093_));
 AOI21_X1 _5290_ (.A(_1093_),
    .B1(_0952_),
    .B2(_0905_),
    .ZN(_1094_));
 XNOR2_X1 _5291_ (.A(_1091_),
    .B(_1094_),
    .ZN(_1095_));
 XNOR2_X1 _5292_ (.A(\fir.p4[11] ),
    .B(_1095_),
    .ZN(_1096_));
 XOR2_X1 _5293_ (.A(_1047_),
    .B(_1096_),
    .Z(_1097_));
 XOR2_X1 _5294_ (.A(\fir.p4[10] ),
    .B(_1097_),
    .Z(_1098_));
 XNOR2_X1 _5295_ (.A(_1045_),
    .B(_1098_),
    .ZN(_1099_));
 XNOR2_X1 _5296_ (.A(_1042_),
    .B(_1099_),
    .ZN(_1100_));
 XNOR2_X1 _5297_ (.A(_1038_),
    .B(_1100_),
    .ZN(_1101_));
 XNOR2_X1 _5298_ (.A(_1036_),
    .B(_1101_),
    .ZN(_1102_));
 XOR2_X1 _5299_ (.A(_1030_),
    .B(_1102_),
    .Z(_1103_));
 XOR2_X1 _5300_ (.A(_1026_),
    .B(_1103_),
    .Z(_1104_));
 XOR2_X1 _5301_ (.A(_1014_),
    .B(_1104_),
    .Z(_1105_));
 XNOR2_X1 _5302_ (.A(_1011_),
    .B(_1105_),
    .ZN(_1106_));
 XOR2_X1 _5303_ (.A(_1009_),
    .B(_1106_),
    .Z(_1107_));
 NAND2_X1 _5304_ (.A1(_0851_),
    .A2(_0964_),
    .ZN(_1108_));
 OAI211_X1 _5305_ (.A(_0966_),
    .B(_0692_),
    .C1(_0851_),
    .C2(_0964_),
    .ZN(_1109_));
 NAND2_X1 _5306_ (.A1(_1108_),
    .A2(_1109_),
    .ZN(_1110_));
 OR2_X1 _5307_ (.A1(_0439_),
    .A2(_0554_),
    .ZN(_1111_));
 AND2_X1 _5308_ (.A1(_0439_),
    .A2(_0554_),
    .ZN(_1112_));
 NOR2_X1 _5309_ (.A1(_0304_),
    .A2(_0416_),
    .ZN(_1113_));
 INV_X1 _5310_ (.A(_0283_),
    .ZN(_1114_));
 INV_X1 _5311_ (.A(_3622_),
    .ZN(_1115_));
 XNOR2_X1 _5312_ (.A(_1115_),
    .B(_0280_),
    .ZN(_1116_));
 AOI22_X1 _5313_ (.A1(_0287_),
    .A2(_3618_),
    .B1(_1115_),
    .B2(_0280_),
    .ZN(_1117_));
 NOR2_X1 _5314_ (.A1(_1115_),
    .A2(_0280_),
    .ZN(_1118_));
 OAI22_X1 _5315_ (.A1(_1114_),
    .A2(_1116_),
    .B1(_1117_),
    .B2(_1118_),
    .ZN(_1119_));
 AOI21_X1 _5316_ (.A(_1113_),
    .B1(_0417_),
    .B2(_1119_),
    .ZN(_1120_));
 OAI21_X1 _5317_ (.A(_1111_),
    .B1(_1112_),
    .B2(_1120_),
    .ZN(_1121_));
 AND3_X1 _5318_ (.A1(_1121_),
    .A2(_0693_),
    .A3(_0965_),
    .ZN(_1122_));
 OAI21_X1 _5319_ (.A(_1107_),
    .B1(_1110_),
    .B2(_1122_),
    .ZN(_1123_));
 NAND3_X1 _5320_ (.A1(_1121_),
    .A2(_0693_),
    .A3(_0965_),
    .ZN(_1124_));
 AND2_X1 _5321_ (.A1(_1108_),
    .A2(_1109_),
    .ZN(_1125_));
 XNOR2_X1 _5322_ (.A(_1009_),
    .B(_1106_),
    .ZN(_1126_));
 NAND3_X1 _5323_ (.A1(_1124_),
    .A2(_1125_),
    .A3(_1126_),
    .ZN(_1127_));
 AOI21_X1 _5324_ (.A(_0575_),
    .B1(_1123_),
    .B2(_1127_),
    .ZN(_1128_));
 AOI21_X1 _5325_ (.A(_1126_),
    .B1(_1125_),
    .B2(_1124_),
    .ZN(_1129_));
 NOR3_X1 _5326_ (.A1(_1122_),
    .A2(_1110_),
    .A3(_1107_),
    .ZN(_1130_));
 NOR3_X1 _5327_ (.A1(\fir.p5[11] ),
    .A2(_1129_),
    .A3(_1130_),
    .ZN(_1131_));
 OAI21_X1 _5328_ (.A(_1007_),
    .B1(_1128_),
    .B2(_1131_),
    .ZN(_1132_));
 OR2_X1 _5329_ (.A1(_0029_),
    .A2(_0970_),
    .ZN(_1133_));
 OAI21_X1 _5330_ (.A(\fir.p5[11] ),
    .B1(_1129_),
    .B2(_1130_),
    .ZN(_1134_));
 NAND3_X1 _5331_ (.A1(_0575_),
    .A2(_1123_),
    .A3(_1127_),
    .ZN(_1135_));
 NAND3_X1 _5332_ (.A1(_1133_),
    .A2(_1134_),
    .A3(_1135_),
    .ZN(_1136_));
 NAND3_X1 _5333_ (.A1(_1006_),
    .A2(_1132_),
    .A3(_1136_),
    .ZN(_1137_));
 XNOR2_X1 _5334_ (.A(\fir.p5[9] ),
    .B(\fir.p5[11] ),
    .ZN(_1138_));
 AOI21_X1 _5335_ (.A(_1133_),
    .B1(_1134_),
    .B2(_1135_),
    .ZN(_1139_));
 NOR3_X1 _5336_ (.A1(_1007_),
    .A2(_1128_),
    .A3(_1131_),
    .ZN(_1140_));
 OAI21_X1 _5337_ (.A(_1138_),
    .B1(_1139_),
    .B2(_1140_),
    .ZN(_1141_));
 NAND3_X1 _5338_ (.A1(_1005_),
    .A2(_1137_),
    .A3(_1141_),
    .ZN(_1142_));
 AND2_X1 _5339_ (.A1(_0849_),
    .A2(_0971_),
    .ZN(_1143_));
 INV_X1 _5340_ (.A(_0847_),
    .ZN(_1144_));
 AOI21_X1 _5341_ (.A(_1143_),
    .B1(_0972_),
    .B2(_1144_),
    .ZN(_1145_));
 NOR3_X1 _5342_ (.A1(_1138_),
    .A2(_1139_),
    .A3(_1140_),
    .ZN(_1146_));
 AOI21_X1 _5343_ (.A(_1006_),
    .B1(_1132_),
    .B2(_1136_),
    .ZN(_1147_));
 OAI21_X1 _5344_ (.A(_1145_),
    .B1(_1146_),
    .B2(_1147_),
    .ZN(_1148_));
 NAND3_X1 _5345_ (.A1(_1002_),
    .A2(_1142_),
    .A3(_1148_),
    .ZN(_1149_));
 XNOR2_X1 _5346_ (.A(_0033_),
    .B(_1001_),
    .ZN(_1150_));
 NOR3_X1 _5347_ (.A1(_1145_),
    .A2(_1146_),
    .A3(_1147_),
    .ZN(_1151_));
 AOI21_X1 _5348_ (.A(_1005_),
    .B1(_1137_),
    .B2(_1141_),
    .ZN(_1152_));
 OAI21_X1 _5349_ (.A(_1150_),
    .B1(_1151_),
    .B2(_1152_),
    .ZN(_1153_));
 NAND3_X1 _5350_ (.A1(_1000_),
    .A2(_1149_),
    .A3(_1153_),
    .ZN(_1154_));
 AND2_X1 _5351_ (.A1(_0846_),
    .A2(_0973_),
    .ZN(_1155_));
 AOI21_X1 _5352_ (.A(_1155_),
    .B1(_0974_),
    .B2(_0844_),
    .ZN(_1156_));
 NOR3_X1 _5353_ (.A1(_1150_),
    .A2(_1151_),
    .A3(_1152_),
    .ZN(_1157_));
 AOI21_X1 _5354_ (.A(_1002_),
    .B1(_1142_),
    .B2(_1148_),
    .ZN(_1158_));
 OAI21_X1 _5355_ (.A(_1156_),
    .B1(_1157_),
    .B2(_1158_),
    .ZN(_1159_));
 NAND3_X1 _5356_ (.A1(_0996_),
    .A2(_1154_),
    .A3(_1159_),
    .ZN(_1160_));
 NOR3_X1 _5357_ (.A1(_1156_),
    .A2(_1157_),
    .A3(_1158_),
    .ZN(_1161_));
 AOI21_X1 _5358_ (.A(_1000_),
    .B1(_1149_),
    .B2(_1153_),
    .ZN(_1162_));
 OAI22_X1 _5359_ (.A1(_0030_),
    .A2(_0843_),
    .B1(_1161_),
    .B2(_1162_),
    .ZN(_1163_));
 NAND3_X1 _5360_ (.A1(_0995_),
    .A2(_1160_),
    .A3(_1163_),
    .ZN(_1164_));
 AND3_X1 _5361_ (.A1(_0996_),
    .A2(_1154_),
    .A3(_1159_),
    .ZN(_1165_));
 AOI21_X1 _5362_ (.A(_0996_),
    .B1(_1154_),
    .B2(_1159_),
    .ZN(_1166_));
 OAI221_X1 _5363_ (.A(_0993_),
    .B1(_1165_),
    .B2(_1166_),
    .C1(_0994_),
    .C2(_0840_),
    .ZN(_1167_));
 NAND2_X1 _5364_ (.A1(_1164_),
    .A2(_1167_),
    .ZN(_1168_));
 NOR2_X1 _5365_ (.A1(_0839_),
    .A2(_0977_),
    .ZN(_1169_));
 AOI21_X1 _5366_ (.A(_1169_),
    .B1(_0978_),
    .B2(_0837_),
    .ZN(_1170_));
 XOR2_X1 _5367_ (.A(_1168_),
    .B(_1170_),
    .Z(_1171_));
 XNOR2_X1 _5368_ (.A(_0984_),
    .B(_1171_),
    .ZN(_1172_));
 XOR2_X1 _5369_ (.A(_0992_),
    .B(_1172_),
    .Z(_1173_));
 XNOR2_X1 _5370_ (.A(_0990_),
    .B(_1173_),
    .ZN(_1174_));
 NOR2_X1 _5371_ (.A1(_0989_),
    .A2(_1174_),
    .ZN(_1175_));
 XOR2_X1 _5372_ (.A(_0031_),
    .B(_2973_),
    .Z(_1176_));
 XOR2_X1 _5373_ (.A(_0989_),
    .B(_1174_),
    .Z(_1177_));
 AOI21_X1 _5374_ (.A(_1175_),
    .B1(_1176_),
    .B2(_1177_),
    .ZN(_1178_));
 NAND2_X1 _5375_ (.A1(\fir.p7[11] ),
    .A2(\fir.p7[10] ),
    .ZN(_1179_));
 XOR2_X1 _5376_ (.A(_0031_),
    .B(_1179_),
    .Z(_1180_));
 AOI22_X1 _5377_ (.A1(_0992_),
    .A2(_1172_),
    .B1(_1173_),
    .B2(_0990_),
    .ZN(_1181_));
 NOR2_X1 _5378_ (.A1(_0984_),
    .A2(_1171_),
    .ZN(_1182_));
 AND4_X1 _5379_ (.A1(_0837_),
    .A2(_0978_),
    .A3(_1164_),
    .A4(_1167_),
    .ZN(_1183_));
 AOI21_X1 _5380_ (.A(_0995_),
    .B1(_1160_),
    .B2(_1163_),
    .ZN(_1184_));
 OR2_X1 _5381_ (.A1(_0839_),
    .A2(_0977_),
    .ZN(_1185_));
 OAI21_X1 _5382_ (.A(_1164_),
    .B1(_1184_),
    .B2(_1185_),
    .ZN(_1186_));
 NOR2_X1 _5383_ (.A1(_1183_),
    .A2(_1186_),
    .ZN(_1187_));
 NOR2_X1 _5384_ (.A1(_1161_),
    .A2(_1165_),
    .ZN(_1188_));
 NOR2_X1 _5385_ (.A1(_0033_),
    .A2(_1001_),
    .ZN(_1189_));
 NOR2_X1 _5386_ (.A1(_1151_),
    .A2(_1157_),
    .ZN(_1190_));
 NAND2_X1 _5387_ (.A1(\fir.p5[9] ),
    .A2(\fir.p5[11] ),
    .ZN(_1191_));
 XOR2_X1 _5388_ (.A(_0036_),
    .B(_1191_),
    .Z(_1192_));
 NOR2_X1 _5389_ (.A1(_1139_),
    .A2(_1146_),
    .ZN(_1193_));
 XOR2_X1 _5390_ (.A(\fir.p5[11] ),
    .B(\fir.p5[10] ),
    .Z(_1194_));
 NAND3_X1 _5391_ (.A1(_0848_),
    .A2(_1123_),
    .A3(_1127_),
    .ZN(_1195_));
 NAND2_X1 _5392_ (.A1(_1014_),
    .A2(_1104_),
    .ZN(_1196_));
 NAND2_X1 _5393_ (.A1(_1011_),
    .A2(_1105_),
    .ZN(_1197_));
 NAND2_X1 _5394_ (.A1(_1196_),
    .A2(_1197_),
    .ZN(_1198_));
 OR2_X1 _5395_ (.A1(_1021_),
    .A2(_1024_),
    .ZN(_1199_));
 OAI21_X1 _5396_ (.A(_1199_),
    .B1(_1025_),
    .B2(_0866_),
    .ZN(_1200_));
 NOR2_X1 _5397_ (.A1(_1026_),
    .A2(_1103_),
    .ZN(_1201_));
 INV_X1 _5398_ (.A(_1102_),
    .ZN(_1202_));
 AOI21_X1 _5399_ (.A(_1201_),
    .B1(_1202_),
    .B2(_1030_),
    .ZN(_1203_));
 NAND2_X1 _5400_ (.A1(_1016_),
    .A2(_1020_),
    .ZN(_1204_));
 OR2_X1 _5401_ (.A1(_0467_),
    .A2(_1018_),
    .ZN(_1205_));
 OAI21_X1 _5402_ (.A(_1205_),
    .B1(_1019_),
    .B2(_0451_),
    .ZN(_1206_));
 XOR2_X1 _5403_ (.A(_0590_),
    .B(_0605_),
    .Z(_1207_));
 XNOR2_X1 _5404_ (.A(_1206_),
    .B(_1207_),
    .ZN(_1208_));
 OR2_X1 _5405_ (.A1(_1031_),
    .A2(_1035_),
    .ZN(_1209_));
 NAND2_X1 _5406_ (.A1(_1032_),
    .A2(_1034_),
    .ZN(_1210_));
 AOI21_X1 _5407_ (.A(_1208_),
    .B1(_1209_),
    .B2(_1210_),
    .ZN(_1211_));
 AND3_X1 _5408_ (.A1(_1210_),
    .A2(_1209_),
    .A3(_1208_),
    .ZN(_1212_));
 OR2_X1 _5409_ (.A1(_1211_),
    .A2(_1212_),
    .ZN(_1213_));
 XNOR2_X1 _5410_ (.A(_1204_),
    .B(_1213_),
    .ZN(_1214_));
 NAND2_X1 _5411_ (.A1(_1038_),
    .A2(_1100_),
    .ZN(_1215_));
 OAI21_X1 _5412_ (.A(_1215_),
    .B1(_1101_),
    .B2(_1036_),
    .ZN(_1216_));
 NAND2_X1 _5413_ (.A1(\fir.p3[11] ),
    .A2(\fir.p3[10] ),
    .ZN(_1217_));
 NOR2_X1 _5414_ (.A1(_0486_),
    .A2(_1040_),
    .ZN(_1218_));
 NOR2_X1 _5415_ (.A1(_0478_),
    .A2(_1041_),
    .ZN(_1219_));
 NOR2_X1 _5416_ (.A1(_1218_),
    .A2(_1219_),
    .ZN(_1220_));
 XNOR2_X1 _5417_ (.A(_1217_),
    .B(_1220_),
    .ZN(_1221_));
 NOR2_X1 _5418_ (.A1(_1045_),
    .A2(_1098_),
    .ZN(_1222_));
 INV_X1 _5419_ (.A(_1099_),
    .ZN(_1223_));
 AOI21_X1 _5420_ (.A(_1222_),
    .B1(_1223_),
    .B2(_1042_),
    .ZN(_1224_));
 XNOR2_X1 _5421_ (.A(_0488_),
    .B(_0624_),
    .ZN(_1225_));
 XNOR2_X1 _5422_ (.A(_0615_),
    .B(_1225_),
    .ZN(_1226_));
 AND3_X1 _5423_ (.A1(_1046_),
    .A2(_0953_),
    .A3(_1096_),
    .ZN(_1227_));
 INV_X1 _5424_ (.A(_1097_),
    .ZN(_1228_));
 AOI21_X1 _5425_ (.A(_1227_),
    .B1(_1228_),
    .B2(\fir.p4[10] ),
    .ZN(_1229_));
 OR2_X1 _5426_ (.A1(_0488_),
    .A2(_1095_),
    .ZN(_1230_));
 NAND2_X1 _5427_ (.A1(_1049_),
    .A2(_1090_),
    .ZN(_1231_));
 OAI211_X1 _5428_ (.A(_1092_),
    .B(_0951_),
    .C1(_1049_),
    .C2(_1090_),
    .ZN(_1232_));
 NAND2_X1 _5429_ (.A1(_0905_),
    .A2(_0952_),
    .ZN(_1233_));
 OAI211_X1 _5430_ (.A(_1231_),
    .B(_1232_),
    .C1(_1091_),
    .C2(_1233_),
    .ZN(_1234_));
 NOR2_X1 _5431_ (.A1(_1052_),
    .A2(_1088_),
    .ZN(_1235_));
 AOI21_X1 _5432_ (.A(_1235_),
    .B1(_1089_),
    .B2(_1050_),
    .ZN(_1236_));
 NOR2_X1 _5433_ (.A1(_0018_),
    .A2(_1053_),
    .ZN(_1237_));
 AND2_X1 _5434_ (.A1(_1056_),
    .A2(_1086_),
    .ZN(_1238_));
 AOI21_X1 _5435_ (.A(_1238_),
    .B1(_1087_),
    .B2(_1054_),
    .ZN(_1239_));
 NAND2_X1 _5436_ (.A1(\fir.p2[9] ),
    .A2(\fir.p2[11] ),
    .ZN(_1240_));
 XOR2_X1 _5437_ (.A(_0024_),
    .B(_1240_),
    .Z(_1241_));
 INV_X1 _5438_ (.A(_1058_),
    .ZN(_1242_));
 NOR2_X1 _5439_ (.A1(_1242_),
    .A2(_1084_),
    .ZN(_1243_));
 AND2_X1 _5440_ (.A1(_1057_),
    .A2(_1085_),
    .ZN(_1244_));
 NOR2_X1 _5441_ (.A1(_1243_),
    .A2(_1244_),
    .ZN(_1245_));
 XOR2_X1 _5442_ (.A(\fir.p2[11] ),
    .B(\fir.p2[10] ),
    .Z(_1246_));
 NAND2_X1 _5443_ (.A1(\fir.p2[11] ),
    .A2(_1083_),
    .ZN(_1247_));
 INV_X1 _5444_ (.A(net286),
    .ZN(_1248_));
 NAND2_X1 _5445_ (.A1(_0937_),
    .A2(_1075_),
    .ZN(_1249_));
 NOR2_X1 _5446_ (.A1(_1060_),
    .A2(_1070_),
    .ZN(_1250_));
 NAND2_X1 _5447_ (.A1(\fir.p1[8] ),
    .A2(_1069_),
    .ZN(_1251_));
 NAND2_X1 _5448_ (.A1(_1067_),
    .A2(_1251_),
    .ZN(_1252_));
 XOR2_X1 _5449_ (.A(_0035_),
    .B(_0924_),
    .Z(_1253_));
 XNOR2_X1 _5450_ (.A(_1062_),
    .B(_1253_),
    .ZN(_1254_));
 XNOR2_X1 _5451_ (.A(\fir.p1[9] ),
    .B(_1254_),
    .ZN(_1255_));
 XNOR2_X1 _5452_ (.A(_1252_),
    .B(_1255_),
    .ZN(_1256_));
 XNOR2_X1 _5453_ (.A(_1250_),
    .B(_1256_),
    .ZN(_1257_));
 XNOR2_X1 _5454_ (.A(_1073_),
    .B(_1257_),
    .ZN(_1258_));
 AND3_X1 _5455_ (.A1(_1249_),
    .A2(_1081_),
    .A3(_1258_),
    .ZN(_1259_));
 AOI21_X1 _5456_ (.A(_1258_),
    .B1(_1081_),
    .B2(_1249_),
    .ZN(_1260_));
 OR2_X1 _5457_ (.A1(_1259_),
    .A2(_1260_),
    .ZN(_1261_));
 XNOR2_X1 _5458_ (.A(_1248_),
    .B(_1261_),
    .ZN(_1262_));
 XNOR2_X1 _5459_ (.A(_1247_),
    .B(_1262_),
    .ZN(_1263_));
 XNOR2_X1 _5460_ (.A(_1246_),
    .B(_1263_),
    .ZN(_1264_));
 XNOR2_X1 _5461_ (.A(_1245_),
    .B(_1264_),
    .ZN(_1265_));
 XNOR2_X1 _5462_ (.A(_1241_),
    .B(_1265_),
    .ZN(_1266_));
 XOR2_X1 _5463_ (.A(_1239_),
    .B(_1266_),
    .Z(_1267_));
 XOR2_X1 _5464_ (.A(_1237_),
    .B(_1267_),
    .Z(_1268_));
 XNOR2_X1 _5465_ (.A(_1236_),
    .B(_1268_),
    .ZN(_1269_));
 XOR2_X1 _5466_ (.A(_1234_),
    .B(_1269_),
    .Z(_1270_));
 XOR2_X1 _5467_ (.A(_1230_),
    .B(_1270_),
    .Z(_1271_));
 XNOR2_X1 _5468_ (.A(_1229_),
    .B(_1271_),
    .ZN(_1272_));
 XOR2_X1 _5469_ (.A(_1226_),
    .B(_1272_),
    .Z(_1273_));
 XNOR2_X1 _5470_ (.A(_1224_),
    .B(_1273_),
    .ZN(_1274_));
 XNOR2_X1 _5471_ (.A(_1221_),
    .B(_1274_),
    .ZN(_1275_));
 XNOR2_X1 _5472_ (.A(_1216_),
    .B(_1275_),
    .ZN(_1276_));
 XNOR2_X1 _5473_ (.A(_1214_),
    .B(_1276_),
    .ZN(_1277_));
 XNOR2_X1 _5474_ (.A(_1203_),
    .B(_1277_),
    .ZN(_1278_));
 XNOR2_X1 _5475_ (.A(_1200_),
    .B(_1278_),
    .ZN(_1279_));
 XOR2_X1 _5476_ (.A(_1198_),
    .B(_1279_),
    .Z(_1280_));
 OR2_X1 _5477_ (.A1(_1009_),
    .A2(_1106_),
    .ZN(_1281_));
 INV_X1 _5478_ (.A(_1281_),
    .ZN(_1282_));
 OAI21_X1 _5479_ (.A(_1280_),
    .B1(_1129_),
    .B2(_1282_),
    .ZN(_1283_));
 OR3_X1 _5480_ (.A1(_1282_),
    .A2(_1129_),
    .A3(_1280_),
    .ZN(_1284_));
 AND3_X1 _5481_ (.A1(\fir.p5[11] ),
    .A2(_1283_),
    .A3(_1284_),
    .ZN(_1285_));
 AOI21_X1 _5482_ (.A(\fir.p5[11] ),
    .B1(_1283_),
    .B2(_1284_),
    .ZN(_1286_));
 OR3_X1 _5483_ (.A1(_1195_),
    .A2(_1285_),
    .A3(_1286_),
    .ZN(_1287_));
 OAI21_X1 _5484_ (.A(_1195_),
    .B1(_1285_),
    .B2(_1286_),
    .ZN(_1288_));
 AND3_X1 _5485_ (.A1(_1194_),
    .A2(_1287_),
    .A3(_1288_),
    .ZN(_1289_));
 AOI21_X1 _5486_ (.A(_1194_),
    .B1(_1287_),
    .B2(_1288_),
    .ZN(_1290_));
 OR3_X1 _5487_ (.A1(_1193_),
    .A2(_1289_),
    .A3(_1290_),
    .ZN(_1291_));
 OAI21_X1 _5488_ (.A(_1193_),
    .B1(_1289_),
    .B2(_1290_),
    .ZN(_1292_));
 AND3_X1 _5489_ (.A1(_1192_),
    .A2(_1291_),
    .A3(_1292_),
    .ZN(_1293_));
 AOI21_X1 _5490_ (.A(_1192_),
    .B1(_1291_),
    .B2(_1292_),
    .ZN(_1294_));
 OR3_X1 _5491_ (.A1(_1190_),
    .A2(_1293_),
    .A3(_1294_),
    .ZN(_1295_));
 OAI21_X1 _5492_ (.A(_1190_),
    .B1(_1293_),
    .B2(_1294_),
    .ZN(_1296_));
 AND3_X1 _5493_ (.A1(_1189_),
    .A2(_1295_),
    .A3(_1296_),
    .ZN(_1297_));
 AOI21_X1 _5494_ (.A(_1189_),
    .B1(_1295_),
    .B2(_1296_),
    .ZN(_1298_));
 OR3_X1 _5495_ (.A1(_1188_),
    .A2(_1297_),
    .A3(_1298_),
    .ZN(_1299_));
 OAI21_X1 _5496_ (.A(_1188_),
    .B1(_1297_),
    .B2(_1298_),
    .ZN(_1300_));
 AND2_X1 _5497_ (.A1(_1299_),
    .A2(_1300_),
    .ZN(_1301_));
 XNOR2_X1 _5498_ (.A(_1187_),
    .B(_1301_),
    .ZN(_1302_));
 XNOR2_X1 _5499_ (.A(_1182_),
    .B(_1302_),
    .ZN(_1303_));
 XOR2_X1 _5500_ (.A(_1181_),
    .B(_1303_),
    .Z(_1304_));
 XNOR2_X1 _5501_ (.A(_1180_),
    .B(_1304_),
    .ZN(_1305_));
 NOR2_X1 _5502_ (.A1(_1178_),
    .A2(_1305_),
    .ZN(_1306_));
 NOR2_X1 _5503_ (.A1(_0031_),
    .A2(_2973_),
    .ZN(_1307_));
 XNOR2_X1 _5504_ (.A(_0037_),
    .B(_1307_),
    .ZN(_1308_));
 XOR2_X1 _5505_ (.A(_1178_),
    .B(_1305_),
    .Z(_1309_));
 AOI21_X1 _5506_ (.A(_1306_),
    .B1(_1308_),
    .B2(_1309_),
    .ZN(_1310_));
 NOR2_X1 _5507_ (.A1(_0031_),
    .A2(_1179_),
    .ZN(_1311_));
 XOR2_X1 _5508_ (.A(_0039_),
    .B(_1311_),
    .Z(_1312_));
 NOR2_X1 _5509_ (.A1(_1181_),
    .A2(_1303_),
    .ZN(_1313_));
 AOI21_X1 _5510_ (.A(_1313_),
    .B1(_1304_),
    .B2(_1180_),
    .ZN(_1314_));
 XNOR2_X1 _5511_ (.A(\fir.p6[11] ),
    .B(\fir.p7[11] ),
    .ZN(_1315_));
 NOR3_X1 _5512_ (.A1(_0984_),
    .A2(_1171_),
    .A3(_1302_),
    .ZN(_1316_));
 OAI211_X1 _5513_ (.A(_1299_),
    .B(_1300_),
    .C1(_1183_),
    .C2(_1186_),
    .ZN(_1317_));
 NAND2_X1 _5514_ (.A1(_1299_),
    .A2(_1317_),
    .ZN(_1318_));
 NAND3_X1 _5515_ (.A1(_1189_),
    .A2(_1295_),
    .A3(_1296_),
    .ZN(_1319_));
 NAND2_X1 _5516_ (.A1(_1295_),
    .A2(_1319_),
    .ZN(_1320_));
 OR2_X1 _5517_ (.A1(_0036_),
    .A2(_1191_),
    .ZN(_1321_));
 NAND3_X1 _5518_ (.A1(_1192_),
    .A2(_1291_),
    .A3(_1292_),
    .ZN(_1322_));
 NAND2_X1 _5519_ (.A1(_1291_),
    .A2(_1322_),
    .ZN(_1323_));
 NAND2_X1 _5520_ (.A1(\fir.p5[11] ),
    .A2(\fir.p5[10] ),
    .ZN(_1324_));
 XNOR2_X1 _5521_ (.A(_0432_),
    .B(_1324_),
    .ZN(_1325_));
 NOR3_X1 _5522_ (.A1(_1195_),
    .A2(_1285_),
    .A3(_1286_),
    .ZN(_1326_));
 AOI21_X1 _5523_ (.A(_1326_),
    .B1(_1288_),
    .B2(_1194_),
    .ZN(_1327_));
 NAND2_X1 _5524_ (.A1(_1283_),
    .A2(_1284_),
    .ZN(_1328_));
 NAND2_X1 _5525_ (.A1(\fir.p5[11] ),
    .A2(_1328_),
    .ZN(_1329_));
 NAND2_X1 _5526_ (.A1(_1198_),
    .A2(_1279_),
    .ZN(_1330_));
 AND2_X1 _5527_ (.A1(_1330_),
    .A2(_1283_),
    .ZN(_1331_));
 INV_X1 _5528_ (.A(_1278_),
    .ZN(_1332_));
 NAND2_X1 _5529_ (.A1(_1200_),
    .A2(_1332_),
    .ZN(_1333_));
 OAI21_X1 _5530_ (.A(_1333_),
    .B1(_1277_),
    .B2(_1203_),
    .ZN(_1334_));
 NOR2_X1 _5531_ (.A1(_1204_),
    .A2(_1213_),
    .ZN(_1335_));
 NOR2_X1 _5532_ (.A1(_1211_),
    .A2(_1335_),
    .ZN(_1336_));
 NOR2_X1 _5533_ (.A1(_1214_),
    .A2(_1276_),
    .ZN(_1337_));
 AOI21_X1 _5534_ (.A(_1337_),
    .B1(_1275_),
    .B2(_1216_),
    .ZN(_1338_));
 AND2_X1 _5535_ (.A1(_1206_),
    .A2(_1207_),
    .ZN(_1339_));
 OR2_X1 _5536_ (.A1(_1217_),
    .A2(_1220_),
    .ZN(_1340_));
 OAI21_X1 _5537_ (.A(_0878_),
    .B1(_0605_),
    .B2(_0590_),
    .ZN(_1341_));
 OAI21_X1 _5538_ (.A(_0859_),
    .B1(\fir.p3[10] ),
    .B2(\fir.p3[9] ),
    .ZN(_1342_));
 XOR2_X1 _5539_ (.A(_1341_),
    .B(_1342_),
    .Z(_1343_));
 XOR2_X1 _5540_ (.A(_1340_),
    .B(_1343_),
    .Z(_1344_));
 XOR2_X1 _5541_ (.A(_1339_),
    .B(_1344_),
    .Z(_1345_));
 INV_X1 _5542_ (.A(_1274_),
    .ZN(_1346_));
 NOR2_X1 _5543_ (.A1(_1221_),
    .A2(_1346_),
    .ZN(_1347_));
 INV_X1 _5544_ (.A(_1224_),
    .ZN(_1348_));
 AOI21_X1 _5545_ (.A(_1347_),
    .B1(_1273_),
    .B2(_1348_),
    .ZN(_1349_));
 OAI22_X1 _5546_ (.A1(_0026_),
    .A2(_0624_),
    .B1(_1225_),
    .B2(_0615_),
    .ZN(_1350_));
 XNOR2_X1 _5547_ (.A(_0465_),
    .B(_1350_),
    .ZN(_1351_));
 OR2_X1 _5548_ (.A1(_1229_),
    .A2(_1271_),
    .ZN(_1352_));
 OAI21_X1 _5549_ (.A(_1352_),
    .B1(_1272_),
    .B2(_1226_),
    .ZN(_1353_));
 NAND2_X1 _5550_ (.A1(_0621_),
    .A2(_0887_),
    .ZN(_1354_));
 MUX2_X1 _5551_ (.A(_0026_),
    .B(_1230_),
    .S(_1270_),
    .Z(_1355_));
 INV_X1 _5552_ (.A(_1355_),
    .ZN(_1356_));
 NAND2_X1 _5553_ (.A1(\fir.p4[11] ),
    .A2(_1270_),
    .ZN(_1357_));
 INV_X1 _5554_ (.A(_1268_),
    .ZN(_1358_));
 NOR2_X1 _5555_ (.A1(_1236_),
    .A2(_1358_),
    .ZN(_1359_));
 AND2_X1 _5556_ (.A1(_1234_),
    .A2(_1269_),
    .ZN(_1360_));
 NOR2_X1 _5557_ (.A1(_1359_),
    .A2(_1360_),
    .ZN(_1361_));
 NOR2_X1 _5558_ (.A1(_1239_),
    .A2(_1266_),
    .ZN(_1362_));
 AOI21_X1 _5559_ (.A(_1362_),
    .B1(_1267_),
    .B2(_1237_),
    .ZN(_1363_));
 NOR2_X1 _5560_ (.A1(_0024_),
    .A2(_1240_),
    .ZN(_1364_));
 OAI21_X1 _5561_ (.A(_1264_),
    .B1(_1244_),
    .B2(_1243_),
    .ZN(_1365_));
 NAND2_X1 _5562_ (.A1(_1241_),
    .A2(_1265_),
    .ZN(_1366_));
 NAND2_X1 _5563_ (.A1(_1365_),
    .A2(_1366_),
    .ZN(_1367_));
 NAND2_X1 _5564_ (.A1(\fir.p2[11] ),
    .A2(\fir.p2[10] ),
    .ZN(_1368_));
 XOR2_X1 _5565_ (.A(_0038_),
    .B(_1368_),
    .Z(_1369_));
 INV_X1 _5566_ (.A(_1263_),
    .ZN(_1370_));
 NAND2_X1 _5567_ (.A1(_1246_),
    .A2(_1370_),
    .ZN(_1371_));
 OAI21_X1 _5568_ (.A(_1371_),
    .B1(_1262_),
    .B2(_1247_),
    .ZN(_1372_));
 NAND2_X1 _5569_ (.A1(\fir.p2[11] ),
    .A2(_1261_),
    .ZN(_1373_));
 INV_X1 _5570_ (.A(_1260_),
    .ZN(_1374_));
 OAI21_X1 _5571_ (.A(_1374_),
    .B1(_1257_),
    .B2(_1073_),
    .ZN(_1375_));
 NAND2_X1 _5572_ (.A1(_1250_),
    .A2(_1256_),
    .ZN(_1376_));
 INV_X1 _5573_ (.A(_1255_),
    .ZN(_1377_));
 NAND2_X1 _5574_ (.A1(_1252_),
    .A2(_1377_),
    .ZN(_1378_));
 INV_X1 _5575_ (.A(_1253_),
    .ZN(_1379_));
 NOR2_X1 _5576_ (.A1(_1062_),
    .A2(_1379_),
    .ZN(_1380_));
 AND2_X1 _5577_ (.A1(\fir.p1[9] ),
    .A2(_1254_),
    .ZN(_1381_));
 NOR2_X1 _5578_ (.A1(_1380_),
    .A2(_1381_),
    .ZN(_1382_));
 OAI21_X1 _5579_ (.A(\fir.p0[11] ),
    .B1(_0035_),
    .B2(_0924_),
    .ZN(_1383_));
 XNOR2_X1 _5580_ (.A(\fir.p1[11] ),
    .B(_1383_),
    .ZN(_1384_));
 XOR2_X1 _5581_ (.A(\fir.p1[10] ),
    .B(_1384_),
    .Z(_1385_));
 XOR2_X1 _5582_ (.A(_1382_),
    .B(_1385_),
    .Z(_1386_));
 XNOR2_X1 _5583_ (.A(_1378_),
    .B(_1386_),
    .ZN(_1387_));
 XOR2_X1 _5584_ (.A(_1376_),
    .B(_1387_),
    .Z(_1388_));
 XNOR2_X1 _5585_ (.A(_1375_),
    .B(_1388_),
    .ZN(_1389_));
 XOR2_X1 _5586_ (.A(_1373_),
    .B(_1389_),
    .Z(_1390_));
 XOR2_X1 _5587_ (.A(_1372_),
    .B(_1390_),
    .Z(_1391_));
 XNOR2_X1 _5588_ (.A(_1369_),
    .B(_1391_),
    .ZN(_1392_));
 XNOR2_X1 _5589_ (.A(_1367_),
    .B(_1392_),
    .ZN(_1393_));
 XOR2_X1 _5590_ (.A(_1364_),
    .B(_1393_),
    .Z(_1394_));
 XNOR2_X1 _5591_ (.A(_1363_),
    .B(_1394_),
    .ZN(_1395_));
 XNOR2_X1 _5592_ (.A(_1361_),
    .B(_1395_),
    .ZN(_1396_));
 XNOR2_X1 _5593_ (.A(_1357_),
    .B(_1396_),
    .ZN(_1397_));
 XNOR2_X1 _5594_ (.A(_1356_),
    .B(_1397_),
    .ZN(_1398_));
 XNOR2_X1 _5595_ (.A(_1354_),
    .B(_1398_),
    .ZN(_1399_));
 INV_X1 _5596_ (.A(_1399_),
    .ZN(_1400_));
 XNOR2_X1 _5597_ (.A(_1353_),
    .B(_1400_),
    .ZN(_1401_));
 XOR2_X1 _5598_ (.A(_1351_),
    .B(_1401_),
    .Z(_1402_));
 XOR2_X1 _5599_ (.A(_1349_),
    .B(_1402_),
    .Z(_1403_));
 XNOR2_X1 _5600_ (.A(_1345_),
    .B(_1403_),
    .ZN(_1404_));
 XOR2_X1 _5601_ (.A(_1338_),
    .B(_1404_),
    .Z(_1405_));
 XNOR2_X1 _5602_ (.A(_1336_),
    .B(_1405_),
    .ZN(_1406_));
 XNOR2_X1 _5603_ (.A(_1334_),
    .B(_1406_),
    .ZN(_1407_));
 XOR2_X1 _5604_ (.A(_1331_),
    .B(_1407_),
    .Z(_1408_));
 XNOR2_X1 _5605_ (.A(_1329_),
    .B(_1408_),
    .ZN(_1409_));
 XNOR2_X1 _5606_ (.A(_1327_),
    .B(_1409_),
    .ZN(_1410_));
 XOR2_X1 _5607_ (.A(_1325_),
    .B(_1410_),
    .Z(_1411_));
 XNOR2_X1 _5608_ (.A(_1323_),
    .B(_1411_),
    .ZN(_1412_));
 XOR2_X1 _5609_ (.A(_1321_),
    .B(_1412_),
    .Z(_1413_));
 XNOR2_X1 _5610_ (.A(_1320_),
    .B(_1413_),
    .ZN(_1414_));
 XNOR2_X1 _5611_ (.A(_1318_),
    .B(_1414_),
    .ZN(_1415_));
 XOR2_X1 _5612_ (.A(_1316_),
    .B(_1415_),
    .Z(_1416_));
 XNOR2_X1 _5613_ (.A(_1315_),
    .B(_1416_),
    .ZN(_1417_));
 XNOR2_X1 _5614_ (.A(_1314_),
    .B(_1417_),
    .ZN(_1418_));
 XNOR2_X1 _5615_ (.A(_1312_),
    .B(_1418_),
    .ZN(_1419_));
 XNOR2_X1 _5616_ (.A(_1310_),
    .B(_1419_),
    .ZN(_1420_));
 NAND2_X1 _5617_ (.A1(_2984_),
    .A2(_1420_),
    .ZN(_1421_));
 INV_X1 _5618_ (.A(_1419_),
    .ZN(_1422_));
 OAI21_X1 _5619_ (.A(_1421_),
    .B1(_1422_),
    .B2(_1310_),
    .ZN(_1423_));
 NOR3_X1 _5620_ (.A1(_0039_),
    .A2(_0031_),
    .A3(_1179_),
    .ZN(_1424_));
 INV_X1 _5621_ (.A(_1417_),
    .ZN(_1425_));
 NOR2_X1 _5622_ (.A1(_1314_),
    .A2(_1425_),
    .ZN(_1426_));
 INV_X1 _5623_ (.A(_1312_),
    .ZN(_1427_));
 AOI21_X1 _5624_ (.A(_1426_),
    .B1(_1418_),
    .B2(_1427_),
    .ZN(_1428_));
 NAND2_X1 _5625_ (.A1(\fir.p6[11] ),
    .A2(_0984_),
    .ZN(_1429_));
 NOR2_X1 _5626_ (.A1(_0984_),
    .A2(_1302_),
    .ZN(_1430_));
 NAND2_X1 _5627_ (.A1(_1171_),
    .A2(_1430_),
    .ZN(_1431_));
 INV_X1 _5628_ (.A(_1416_),
    .ZN(_1432_));
 OAI22_X1 _5629_ (.A1(_1431_),
    .A2(_1415_),
    .B1(_1432_),
    .B2(_1315_),
    .ZN(_1433_));
 NAND2_X1 _5630_ (.A1(\fir.p7[11] ),
    .A2(_1302_),
    .ZN(_1434_));
 NOR2_X1 _5631_ (.A1(_1434_),
    .A2(_1415_),
    .ZN(_1435_));
 NAND2_X1 _5632_ (.A1(_1323_),
    .A2(_1411_),
    .ZN(_1436_));
 OAI21_X1 _5633_ (.A(_1436_),
    .B1(_1412_),
    .B2(_1321_),
    .ZN(_1437_));
 NOR2_X1 _5634_ (.A1(_0021_),
    .A2(_1324_),
    .ZN(_1438_));
 OAI21_X1 _5635_ (.A(_1409_),
    .B1(_1289_),
    .B2(_1326_),
    .ZN(_1439_));
 NAND2_X1 _5636_ (.A1(_1325_),
    .A2(_1410_),
    .ZN(_1440_));
 AND2_X1 _5637_ (.A1(_1439_),
    .A2(_1440_),
    .ZN(_1441_));
 XNOR2_X1 _5638_ (.A(\fir.p5[11] ),
    .B(\fir.p5[10] ),
    .ZN(_1442_));
 NOR2_X1 _5639_ (.A1(_1329_),
    .A2(_1408_),
    .ZN(_1443_));
 NAND2_X1 _5640_ (.A1(_1334_),
    .A2(_1406_),
    .ZN(_1444_));
 OAI21_X1 _5641_ (.A(_1444_),
    .B1(_1407_),
    .B2(_1331_),
    .ZN(_1445_));
 OR2_X1 _5642_ (.A1(_1338_),
    .A2(_1404_),
    .ZN(_1446_));
 AND2_X1 _5643_ (.A1(_1338_),
    .A2(_1404_),
    .ZN(_1447_));
 OAI21_X1 _5644_ (.A(_1446_),
    .B1(_1447_),
    .B2(_1336_),
    .ZN(_1448_));
 NAND2_X1 _5645_ (.A1(_1339_),
    .A2(_1344_),
    .ZN(_1449_));
 OAI21_X1 _5646_ (.A(_1449_),
    .B1(_1343_),
    .B2(_1340_),
    .ZN(_1450_));
 NOR2_X1 _5647_ (.A1(_1349_),
    .A2(_1402_),
    .ZN(_1451_));
 AOI21_X1 _5648_ (.A(_1451_),
    .B1(_1403_),
    .B2(_1345_),
    .ZN(_1452_));
 OAI211_X1 _5649_ (.A(_0859_),
    .B(_1341_),
    .C1(\fir.p3[9] ),
    .C2(\fir.p3[10] ),
    .ZN(_1453_));
 NAND2_X1 _5650_ (.A1(\fir.p3[11] ),
    .A2(_1350_),
    .ZN(_1454_));
 NAND2_X1 _5651_ (.A1(_0859_),
    .A2(_1031_),
    .ZN(_1455_));
 NOR2_X1 _5652_ (.A1(\fir.p3[11] ),
    .A2(\fir.p3[10] ),
    .ZN(_1456_));
 AOI21_X1 _5653_ (.A(_1456_),
    .B1(_1217_),
    .B2(\fir.p3[9] ),
    .ZN(_1457_));
 XNOR2_X1 _5654_ (.A(_1455_),
    .B(_1457_),
    .ZN(_1458_));
 XOR2_X1 _5655_ (.A(_1454_),
    .B(_1458_),
    .Z(_1459_));
 XNOR2_X1 _5656_ (.A(_1453_),
    .B(_1459_),
    .ZN(_1460_));
 OAI21_X1 _5657_ (.A(_0887_),
    .B1(_0898_),
    .B2(_0026_),
    .ZN(_1461_));
 XNOR2_X1 _5658_ (.A(_0465_),
    .B(_1461_),
    .ZN(_1462_));
 NAND2_X1 _5659_ (.A1(_1356_),
    .A2(_1397_),
    .ZN(_1463_));
 OR2_X1 _5660_ (.A1(_1354_),
    .A2(_1398_),
    .ZN(_1464_));
 NAND2_X1 _5661_ (.A1(_1463_),
    .A2(_1464_),
    .ZN(_1465_));
 NOR2_X1 _5662_ (.A1(\fir.p4[11] ),
    .A2(\fir.p4[10] ),
    .ZN(_1466_));
 AOI21_X1 _5663_ (.A(_1466_),
    .B1(_0896_),
    .B2(\fir.p4[9] ),
    .ZN(_1467_));
 MUX2_X1 _5664_ (.A(_0026_),
    .B(_1357_),
    .S(_1396_),
    .Z(_1468_));
 NAND2_X1 _5665_ (.A1(\fir.p4[11] ),
    .A2(_1396_),
    .ZN(_1469_));
 OAI21_X1 _5666_ (.A(_1395_),
    .B1(_1360_),
    .B2(_1359_),
    .ZN(_1470_));
 INV_X1 _5667_ (.A(_1394_),
    .ZN(_1471_));
 OAI21_X1 _5668_ (.A(_1470_),
    .B1(_1471_),
    .B2(_1363_),
    .ZN(_1472_));
 AOI21_X1 _5669_ (.A(_1392_),
    .B1(_1366_),
    .B2(_1365_),
    .ZN(_1473_));
 AOI21_X1 _5670_ (.A(_1473_),
    .B1(_1393_),
    .B2(_1364_),
    .ZN(_1474_));
 NOR2_X1 _5671_ (.A1(_0038_),
    .A2(_1368_),
    .ZN(_1475_));
 AND2_X1 _5672_ (.A1(_1372_),
    .A2(_1390_),
    .ZN(_1476_));
 AOI21_X1 _5673_ (.A(_1476_),
    .B1(_1391_),
    .B2(_1369_),
    .ZN(_1477_));
 NAND3_X1 _5674_ (.A1(\fir.p2[11] ),
    .A2(_1261_),
    .A3(_1389_),
    .ZN(_1478_));
 OR2_X1 _5675_ (.A1(_1376_),
    .A2(_1387_),
    .ZN(_1479_));
 NAND2_X1 _5676_ (.A1(_1375_),
    .A2(_1388_),
    .ZN(_1480_));
 NOR3_X1 _5677_ (.A1(\fir.p1[11] ),
    .A2(_0035_),
    .A3(_0924_),
    .ZN(_1481_));
 AOI21_X1 _5678_ (.A(_1481_),
    .B1(_1384_),
    .B2(\fir.p1[10] ),
    .ZN(_1482_));
 INV_X1 _5679_ (.A(net128),
    .ZN(_1483_));
 NOR2_X1 _5680_ (.A1(\fir.p1[11] ),
    .A2(_1483_),
    .ZN(_1484_));
 XNOR2_X1 _5681_ (.A(_1482_),
    .B(_1484_),
    .ZN(_1485_));
 OAI21_X1 _5682_ (.A(_1385_),
    .B1(_1381_),
    .B2(_1380_),
    .ZN(_1486_));
 OAI21_X1 _5683_ (.A(_1486_),
    .B1(_1386_),
    .B2(_1378_),
    .ZN(_1487_));
 XNOR2_X1 _5684_ (.A(_1485_),
    .B(_1487_),
    .ZN(_1488_));
 AND3_X1 _5685_ (.A1(_1479_),
    .A2(_1480_),
    .A3(_1488_),
    .ZN(_1489_));
 AOI21_X1 _5686_ (.A(_1488_),
    .B1(_1480_),
    .B2(_1479_),
    .ZN(_1490_));
 OR2_X1 _5687_ (.A1(_1489_),
    .A2(_1490_),
    .ZN(_1491_));
 XOR2_X1 _5688_ (.A(_1478_),
    .B(_1491_),
    .Z(_1492_));
 XNOR2_X1 _5689_ (.A(_1246_),
    .B(_1492_),
    .ZN(_1493_));
 XOR2_X1 _5690_ (.A(_1477_),
    .B(_1493_),
    .Z(_1494_));
 XOR2_X1 _5691_ (.A(_1475_),
    .B(_1494_),
    .Z(_1495_));
 XNOR2_X1 _5692_ (.A(_1474_),
    .B(_1495_),
    .ZN(_1496_));
 XOR2_X1 _5693_ (.A(_1472_),
    .B(_1496_),
    .Z(_1497_));
 XOR2_X1 _5694_ (.A(_1469_),
    .B(_1497_),
    .Z(_1498_));
 XNOR2_X1 _5695_ (.A(_1468_),
    .B(_1498_),
    .ZN(_1499_));
 XOR2_X1 _5696_ (.A(_1467_),
    .B(_1499_),
    .Z(_1500_));
 XNOR2_X1 _5697_ (.A(_1465_),
    .B(_1500_),
    .ZN(_1501_));
 XNOR2_X1 _5698_ (.A(_1462_),
    .B(_1501_),
    .ZN(_1502_));
 INV_X1 _5699_ (.A(_1401_),
    .ZN(_1503_));
 NAND2_X1 _5700_ (.A1(_1351_),
    .A2(_1503_),
    .ZN(_1504_));
 NAND2_X1 _5701_ (.A1(_1353_),
    .A2(_1400_),
    .ZN(_1505_));
 AOI21_X1 _5702_ (.A(_1502_),
    .B1(_1504_),
    .B2(_1505_),
    .ZN(_1506_));
 AND3_X1 _5703_ (.A1(_1505_),
    .A2(_1504_),
    .A3(_1502_),
    .ZN(_1507_));
 NOR2_X1 _5704_ (.A1(_1506_),
    .A2(_1507_),
    .ZN(_1508_));
 XNOR2_X1 _5705_ (.A(_1460_),
    .B(_1508_),
    .ZN(_1509_));
 XOR2_X1 _5706_ (.A(_1452_),
    .B(_1509_),
    .Z(_1510_));
 XOR2_X1 _5707_ (.A(_1450_),
    .B(_1510_),
    .Z(_1511_));
 XNOR2_X1 _5708_ (.A(_1448_),
    .B(_1511_),
    .ZN(_1512_));
 XNOR2_X1 _5709_ (.A(_1445_),
    .B(_1512_),
    .ZN(_1513_));
 XNOR2_X1 _5710_ (.A(_1443_),
    .B(_1513_),
    .ZN(_1514_));
 XNOR2_X1 _5711_ (.A(_1442_),
    .B(_1514_),
    .ZN(_1515_));
 XOR2_X1 _5712_ (.A(_1441_),
    .B(_1515_),
    .Z(_1516_));
 XOR2_X1 _5713_ (.A(_1438_),
    .B(_1516_),
    .Z(_1517_));
 XOR2_X1 _5714_ (.A(_1437_),
    .B(_1517_),
    .Z(_1518_));
 AOI21_X1 _5715_ (.A(_1414_),
    .B1(_1317_),
    .B2(_1299_),
    .ZN(_1519_));
 AND2_X1 _5716_ (.A1(_1320_),
    .A2(_1413_),
    .ZN(_1520_));
 OAI21_X1 _5717_ (.A(_1518_),
    .B1(_1519_),
    .B2(_1520_),
    .ZN(_1521_));
 OR3_X1 _5718_ (.A1(_1520_),
    .A2(_1519_),
    .A3(_1518_),
    .ZN(_1522_));
 NAND2_X1 _5719_ (.A1(_1521_),
    .A2(_1522_),
    .ZN(_1523_));
 NOR2_X1 _5720_ (.A1(_0016_),
    .A2(_1415_),
    .ZN(_1524_));
 XNOR2_X1 _5721_ (.A(_1523_),
    .B(_1524_),
    .ZN(_1525_));
 XNOR2_X1 _5722_ (.A(_1435_),
    .B(_1525_),
    .ZN(_1526_));
 XOR2_X1 _5723_ (.A(_1315_),
    .B(_1526_),
    .Z(_1527_));
 XNOR2_X1 _5724_ (.A(_1433_),
    .B(_1527_),
    .ZN(_1528_));
 XNOR2_X1 _5725_ (.A(_1429_),
    .B(_1528_),
    .ZN(_1529_));
 XNOR2_X1 _5726_ (.A(_1428_),
    .B(_1529_),
    .ZN(_1530_));
 XNOR2_X1 _5727_ (.A(_1424_),
    .B(_1530_),
    .ZN(_1531_));
 AND2_X1 _5728_ (.A1(_1423_),
    .A2(_1531_),
    .ZN(_1532_));
 NOR2_X1 _5729_ (.A1(_1428_),
    .A2(_1529_),
    .ZN(_1533_));
 NAND2_X1 _5730_ (.A1(_1428_),
    .A2(_1529_),
    .ZN(_1534_));
 AOI21_X1 _5731_ (.A(_1533_),
    .B1(_1534_),
    .B2(_1424_),
    .ZN(_1535_));
 INV_X1 _5732_ (.A(net169),
    .ZN(_1536_));
 NOR2_X1 _5733_ (.A1(_1536_),
    .A2(_0984_),
    .ZN(_1537_));
 NAND2_X1 _5734_ (.A1(_1433_),
    .A2(_1527_),
    .ZN(_1538_));
 OAI21_X1 _5735_ (.A(_1538_),
    .B1(_1528_),
    .B2(_1429_),
    .ZN(_1539_));
 NAND2_X1 _5736_ (.A1(_1523_),
    .A2(_1524_),
    .ZN(_1540_));
 NAND2_X1 _5737_ (.A1(_1438_),
    .A2(_1516_),
    .ZN(_1541_));
 OAI21_X1 _5738_ (.A(_1541_),
    .B1(_1515_),
    .B2(_1441_),
    .ZN(_1542_));
 NOR2_X1 _5739_ (.A1(_1442_),
    .A2(_1514_),
    .ZN(_1543_));
 INV_X1 _5740_ (.A(_1513_),
    .ZN(_1544_));
 NOR3_X1 _5741_ (.A1(_0575_),
    .A2(_1328_),
    .A3(_1408_),
    .ZN(_1545_));
 AOI21_X1 _5742_ (.A(_1543_),
    .B1(_1544_),
    .B2(_1545_),
    .ZN(_1546_));
 INV_X1 _5743_ (.A(_1546_),
    .ZN(_1547_));
 INV_X1 _5744_ (.A(_1512_),
    .ZN(_1548_));
 AOI22_X1 _5745_ (.A1(_1448_),
    .A2(_1511_),
    .B1(_1548_),
    .B2(_1445_),
    .ZN(_1549_));
 NOR2_X1 _5746_ (.A1(_1452_),
    .A2(_1509_),
    .ZN(_1550_));
 AOI21_X1 _5747_ (.A(_1550_),
    .B1(_1510_),
    .B2(_1450_),
    .ZN(_1551_));
 INV_X1 _5748_ (.A(_1453_),
    .ZN(_1552_));
 NAND2_X1 _5749_ (.A1(_1552_),
    .A2(_1459_),
    .ZN(_1553_));
 OAI21_X1 _5750_ (.A(_1553_),
    .B1(_1458_),
    .B2(_1454_),
    .ZN(_1554_));
 NAND2_X1 _5751_ (.A1(_1455_),
    .A2(_1457_),
    .ZN(_1555_));
 NAND2_X1 _5752_ (.A1(\fir.p3[11] ),
    .A2(_1461_),
    .ZN(_1556_));
 INV_X1 _5753_ (.A(_0858_),
    .ZN(_1557_));
 OAI21_X1 _5754_ (.A(_1017_),
    .B1(_1557_),
    .B2(\fir.p3[11] ),
    .ZN(_1558_));
 XOR2_X1 _5755_ (.A(_1556_),
    .B(_1558_),
    .Z(_1559_));
 XNOR2_X1 _5756_ (.A(_1555_),
    .B(_1559_),
    .ZN(_1560_));
 AOI21_X1 _5757_ (.A(_1500_),
    .B1(_1464_),
    .B2(_1463_),
    .ZN(_1561_));
 AOI21_X1 _5758_ (.A(_1561_),
    .B1(_1501_),
    .B2(_1462_),
    .ZN(_1562_));
 XNOR2_X1 _5759_ (.A(_0465_),
    .B(_1040_),
    .ZN(_1563_));
 NOR2_X1 _5760_ (.A1(_1468_),
    .A2(_1498_),
    .ZN(_1564_));
 NAND2_X1 _5761_ (.A1(_1468_),
    .A2(_1498_),
    .ZN(_1565_));
 AOI21_X1 _5762_ (.A(_1564_),
    .B1(_1565_),
    .B2(_1467_),
    .ZN(_1566_));
 INV_X1 _5763_ (.A(_1495_),
    .ZN(_1567_));
 NOR2_X1 _5764_ (.A1(_1474_),
    .A2(_1567_),
    .ZN(_1568_));
 AOI21_X1 _5765_ (.A(_1568_),
    .B1(_1496_),
    .B2(_1472_),
    .ZN(_1569_));
 NAND2_X1 _5766_ (.A1(_1475_),
    .A2(_1494_),
    .ZN(_1570_));
 OAI21_X1 _5767_ (.A(_1570_),
    .B1(_1493_),
    .B2(_1477_),
    .ZN(_1571_));
 NAND3_X1 _5768_ (.A1(\fir.p2[11] ),
    .A2(_1389_),
    .A3(_1491_),
    .ZN(_1572_));
 AOI21_X1 _5769_ (.A(\fir.p1[11] ),
    .B1(\fir.p0[11] ),
    .B2(_1482_),
    .ZN(_1573_));
 NOR2_X1 _5770_ (.A1(_1378_),
    .A2(_1386_),
    .ZN(_1574_));
 AOI21_X1 _5771_ (.A(_1490_),
    .B1(_1485_),
    .B2(_1574_),
    .ZN(_1575_));
 INV_X1 _5772_ (.A(_1485_),
    .ZN(_1576_));
 OAI21_X1 _5773_ (.A(_1575_),
    .B1(_1576_),
    .B2(_1486_),
    .ZN(_1577_));
 NOR2_X1 _5774_ (.A1(_1573_),
    .A2(_1577_),
    .ZN(_1578_));
 XNOR2_X1 _5775_ (.A(_1572_),
    .B(_1578_),
    .ZN(_1579_));
 AND2_X1 _5776_ (.A1(_1246_),
    .A2(_1492_),
    .ZN(_1580_));
 NOR2_X1 _5777_ (.A1(_1261_),
    .A2(_1572_),
    .ZN(_1581_));
 OAI21_X1 _5778_ (.A(_1579_),
    .B1(_1580_),
    .B2(_1581_),
    .ZN(_1582_));
 OR3_X1 _5779_ (.A1(_1581_),
    .A2(_1580_),
    .A3(_1579_),
    .ZN(_1583_));
 NAND2_X1 _5780_ (.A1(_1582_),
    .A2(_1583_),
    .ZN(_1584_));
 XOR2_X1 _5781_ (.A(_1368_),
    .B(_1584_),
    .Z(_1585_));
 XNOR2_X1 _5782_ (.A(_1571_),
    .B(_1585_),
    .ZN(_1586_));
 XOR2_X1 _5783_ (.A(_1569_),
    .B(_1586_),
    .Z(_1587_));
 NOR2_X1 _5784_ (.A1(_0488_),
    .A2(_1497_),
    .ZN(_1588_));
 XNOR2_X1 _5785_ (.A(_1587_),
    .B(_1588_),
    .ZN(_1589_));
 MUX2_X1 _5786_ (.A(_0026_),
    .B(_1469_),
    .S(_1497_),
    .Z(_1590_));
 XNOR2_X1 _5787_ (.A(\fir.p4[11] ),
    .B(_0026_),
    .ZN(_1591_));
 XNOR2_X1 _5788_ (.A(_1590_),
    .B(_1591_),
    .ZN(_1592_));
 XOR2_X1 _5789_ (.A(_1589_),
    .B(_1592_),
    .Z(_1593_));
 XNOR2_X1 _5790_ (.A(_1566_),
    .B(_1593_),
    .ZN(_1594_));
 XNOR2_X1 _5791_ (.A(_1563_),
    .B(_1594_),
    .ZN(_1595_));
 XOR2_X1 _5792_ (.A(_1562_),
    .B(_1595_),
    .Z(_1596_));
 XOR2_X1 _5793_ (.A(_1560_),
    .B(_1596_),
    .Z(_1597_));
 AND2_X1 _5794_ (.A1(_1460_),
    .A2(_1508_),
    .ZN(_1598_));
 OAI21_X1 _5795_ (.A(_1597_),
    .B1(_1598_),
    .B2(_1506_),
    .ZN(_1599_));
 OR3_X1 _5796_ (.A1(_1506_),
    .A2(_1598_),
    .A3(_1597_),
    .ZN(_1600_));
 AND2_X1 _5797_ (.A1(_1599_),
    .A2(_1600_),
    .ZN(_1601_));
 XNOR2_X1 _5798_ (.A(_1554_),
    .B(_1601_),
    .ZN(_1602_));
 XOR2_X1 _5799_ (.A(_1551_),
    .B(_1602_),
    .Z(_1603_));
 XNOR2_X1 _5800_ (.A(_1549_),
    .B(_1603_),
    .ZN(_1604_));
 XNOR2_X1 _5801_ (.A(_0029_),
    .B(_1604_),
    .ZN(_1605_));
 OAI21_X1 _5802_ (.A(\fir.p5[11] ),
    .B1(_1408_),
    .B2(_1513_),
    .ZN(_1606_));
 XNOR2_X1 _5803_ (.A(_1605_),
    .B(_1606_),
    .ZN(_1607_));
 XNOR2_X1 _5804_ (.A(_1547_),
    .B(_1607_),
    .ZN(_1608_));
 XOR2_X1 _5805_ (.A(_1324_),
    .B(_1608_),
    .Z(_1609_));
 XOR2_X1 _5806_ (.A(_1542_),
    .B(_1609_),
    .Z(_1610_));
 INV_X1 _5807_ (.A(_1610_),
    .ZN(_1611_));
 AND2_X1 _5808_ (.A1(_1437_),
    .A2(_1517_),
    .ZN(_1612_));
 INV_X1 _5809_ (.A(_1612_),
    .ZN(_1613_));
 AOI21_X1 _5810_ (.A(_1611_),
    .B1(_1521_),
    .B2(_1613_),
    .ZN(_1614_));
 AND3_X1 _5811_ (.A1(_1613_),
    .A2(_1521_),
    .A3(_1611_),
    .ZN(_1615_));
 OR2_X1 _5812_ (.A1(_1614_),
    .A2(_1615_),
    .ZN(_1616_));
 XNOR2_X1 _5813_ (.A(_1540_),
    .B(_1616_),
    .ZN(_1617_));
 XOR2_X1 _5814_ (.A(_1315_),
    .B(_1617_),
    .Z(_1618_));
 NOR2_X1 _5815_ (.A1(_1315_),
    .A2(_1526_),
    .ZN(_1619_));
 AND2_X1 _5816_ (.A1(_1435_),
    .A2(_1525_),
    .ZN(_1620_));
 OAI21_X1 _5817_ (.A(_1618_),
    .B1(_1619_),
    .B2(_1620_),
    .ZN(_1621_));
 OR3_X1 _5818_ (.A1(_1620_),
    .A2(_1619_),
    .A3(_1618_),
    .ZN(_1622_));
 AND2_X1 _5819_ (.A1(_1621_),
    .A2(_1622_),
    .ZN(_1623_));
 XNOR2_X1 _5820_ (.A(_1429_),
    .B(_1623_),
    .ZN(_1624_));
 XOR2_X1 _5821_ (.A(_1539_),
    .B(_1624_),
    .Z(_1625_));
 XNOR2_X1 _5822_ (.A(_1537_),
    .B(_1625_),
    .ZN(_1626_));
 XOR2_X1 _5823_ (.A(_1535_),
    .B(_1626_),
    .Z(_1627_));
 XOR2_X1 _5824_ (.A(_1532_),
    .B(_1627_),
    .Z(_1628_));
 XOR2_X1 _5825_ (.A(_2984_),
    .B(_1420_),
    .Z(_1629_));
 NAND2_X1 _5826_ (.A1(\fir.p7[10] ),
    .A2(\fir.p7[8] ),
    .ZN(_1630_));
 NOR3_X1 _5827_ (.A1(_0031_),
    .A2(_0034_),
    .A3(_1630_),
    .ZN(_1631_));
 OR2_X1 _5828_ (.A1(\fir.p7[10] ),
    .A2(\fir.p7[8] ),
    .ZN(_1632_));
 XNOR2_X1 _5829_ (.A(_0724_),
    .B(_0725_),
    .ZN(_1633_));
 XNOR2_X1 _5830_ (.A(_0833_),
    .B(_1633_),
    .ZN(_1634_));
 NOR2_X1 _5831_ (.A1(_0984_),
    .A2(_1634_),
    .ZN(_1635_));
 XOR2_X1 _5832_ (.A(_0981_),
    .B(_1635_),
    .Z(_1636_));
 NAND3_X1 _5833_ (.A1(_1632_),
    .A2(_1630_),
    .A3(_1636_),
    .ZN(_1637_));
 NAND2_X1 _5834_ (.A1(_0985_),
    .A2(_1634_),
    .ZN(_1638_));
 NAND2_X1 _5835_ (.A1(_1637_),
    .A2(_1638_),
    .ZN(_1639_));
 XNOR2_X1 _5836_ (.A(_0988_),
    .B(_0986_),
    .ZN(_1640_));
 AND2_X1 _5837_ (.A1(_1639_),
    .A2(_1640_),
    .ZN(_1641_));
 XOR2_X1 _5838_ (.A(_0031_),
    .B(_1630_),
    .Z(_1642_));
 OR2_X1 _5839_ (.A1(_1639_),
    .A2(_1640_),
    .ZN(_1643_));
 AOI21_X1 _5840_ (.A(_1641_),
    .B1(_1642_),
    .B2(_1643_),
    .ZN(_1644_));
 XNOR2_X1 _5841_ (.A(_1176_),
    .B(_1177_),
    .ZN(_1645_));
 NOR2_X1 _5842_ (.A1(_1644_),
    .A2(_1645_),
    .ZN(_1646_));
 NOR2_X1 _5843_ (.A1(_0031_),
    .A2(_1630_),
    .ZN(_1647_));
 XNOR2_X1 _5844_ (.A(_0034_),
    .B(_1647_),
    .ZN(_1648_));
 XOR2_X1 _5845_ (.A(_1644_),
    .B(_1645_),
    .Z(_1649_));
 AOI21_X1 _5846_ (.A(_1646_),
    .B1(_1648_),
    .B2(_1649_),
    .ZN(_1650_));
 XNOR2_X1 _5847_ (.A(_1308_),
    .B(_1309_),
    .ZN(_1651_));
 XOR2_X1 _5848_ (.A(_1650_),
    .B(_1651_),
    .Z(_1652_));
 AND2_X1 _5849_ (.A1(_1631_),
    .A2(_1652_),
    .ZN(_1653_));
 NOR2_X1 _5850_ (.A1(_1650_),
    .A2(_1651_),
    .ZN(_1654_));
 OAI21_X1 _5851_ (.A(_1629_),
    .B1(_1653_),
    .B2(_1654_),
    .ZN(_1655_));
 XNOR2_X1 _5852_ (.A(_1423_),
    .B(_1531_),
    .ZN(_1656_));
 NOR2_X1 _5853_ (.A1(_1655_),
    .A2(_1656_),
    .ZN(_1657_));
 NAND4_X1 _5854_ (.A1(\fir.p6[11] ),
    .A2(\fir.p6[10] ),
    .A3(\fir.p7[9] ),
    .A4(\fir.p7[7] ),
    .ZN(_1658_));
 XOR2_X1 _5855_ (.A(_0032_),
    .B(_1658_),
    .Z(_1659_));
 AOI22_X1 _5856_ (.A1(\fir.p6[11] ),
    .A2(\fir.p6[10] ),
    .B1(\fir.p7[9] ),
    .B2(\fir.p7[7] ),
    .ZN(_1660_));
 INV_X1 _5857_ (.A(_1660_),
    .ZN(_1661_));
 NAND2_X1 _5858_ (.A1(_1661_),
    .A2(_1658_),
    .ZN(_1662_));
 XOR2_X1 _5859_ (.A(_0747_),
    .B(_0748_),
    .Z(_1663_));
 XNOR2_X1 _5860_ (.A(_1663_),
    .B(_0832_),
    .ZN(_1664_));
 AND2_X1 _5861_ (.A1(\fir.p7[10] ),
    .A2(_1664_),
    .ZN(_1665_));
 INV_X1 _5862_ (.A(_1665_),
    .ZN(_1666_));
 XNOR2_X1 _5863_ (.A(_0991_),
    .B(_1634_),
    .ZN(_1667_));
 NOR2_X1 _5864_ (.A1(_1666_),
    .A2(_1667_),
    .ZN(_1668_));
 XOR2_X1 _5865_ (.A(\fir.p7[9] ),
    .B(\fir.p7[7] ),
    .Z(_1669_));
 XNOR2_X1 _5866_ (.A(_1665_),
    .B(_1667_),
    .ZN(_1670_));
 AOI21_X1 _5867_ (.A(_1668_),
    .B1(_1669_),
    .B2(_1670_),
    .ZN(_1671_));
 NAND2_X1 _5868_ (.A1(_1632_),
    .A2(_1630_),
    .ZN(_1672_));
 XNOR2_X1 _5869_ (.A(_1672_),
    .B(_1636_),
    .ZN(_1673_));
 XOR2_X1 _5870_ (.A(_1671_),
    .B(_1673_),
    .Z(_1674_));
 NOR2_X1 _5871_ (.A1(_1662_),
    .A2(_1674_),
    .ZN(_1675_));
 INV_X1 _5872_ (.A(_1671_),
    .ZN(_1676_));
 AOI21_X1 _5873_ (.A(_1675_),
    .B1(_1673_),
    .B2(_1676_),
    .ZN(_1677_));
 XNOR2_X1 _5874_ (.A(_1639_),
    .B(_1640_),
    .ZN(_1678_));
 XNOR2_X1 _5875_ (.A(_1642_),
    .B(_1678_),
    .ZN(_1679_));
 XNOR2_X1 _5876_ (.A(_1677_),
    .B(_1679_),
    .ZN(_1680_));
 NAND2_X1 _5877_ (.A1(_1659_),
    .A2(_1680_),
    .ZN(_1681_));
 INV_X1 _5878_ (.A(_1679_),
    .ZN(_1682_));
 OAI21_X1 _5879_ (.A(_1681_),
    .B1(_1682_),
    .B2(_1677_),
    .ZN(_1683_));
 XOR2_X1 _5880_ (.A(_1648_),
    .B(_1649_),
    .Z(_1684_));
 NAND2_X1 _5881_ (.A1(_1683_),
    .A2(_1684_),
    .ZN(_1685_));
 NOR2_X1 _5882_ (.A1(_0032_),
    .A2(_1658_),
    .ZN(_1686_));
 XOR2_X1 _5883_ (.A(_1683_),
    .B(_1684_),
    .Z(_1687_));
 NAND2_X1 _5884_ (.A1(_1686_),
    .A2(_1687_),
    .ZN(_1688_));
 NAND2_X1 _5885_ (.A1(_1685_),
    .A2(_1688_),
    .ZN(_1689_));
 XOR2_X1 _5886_ (.A(_1631_),
    .B(_1652_),
    .Z(_1690_));
 AND2_X1 _5887_ (.A1(_1689_),
    .A2(_1690_),
    .ZN(_1691_));
 OR3_X1 _5888_ (.A1(_1654_),
    .A2(_1653_),
    .A3(_1629_),
    .ZN(_1692_));
 AND2_X1 _5889_ (.A1(_1655_),
    .A2(_1692_),
    .ZN(_1693_));
 AND2_X1 _5890_ (.A1(_1691_),
    .A2(_1693_),
    .ZN(_1694_));
 XOR2_X1 _5891_ (.A(_1655_),
    .B(_1656_),
    .Z(_1695_));
 XOR2_X1 _5892_ (.A(_1691_),
    .B(_1693_),
    .Z(_1696_));
 AND2_X1 _5893_ (.A1(_1696_),
    .A2(_1695_),
    .ZN(_1697_));
 XOR2_X1 _5894_ (.A(_1669_),
    .B(_1670_),
    .Z(_1698_));
 XOR2_X1 _5895_ (.A(\fir.p7[8] ),
    .B(\fir.p7[6] ),
    .Z(_1699_));
 XOR2_X1 _5896_ (.A(\fir.p7[10] ),
    .B(_1664_),
    .Z(_1700_));
 XOR2_X1 _5897_ (.A(_0830_),
    .B(_0831_),
    .Z(_1701_));
 AND2_X1 _5898_ (.A1(\fir.p7[9] ),
    .A2(_1701_),
    .ZN(_1702_));
 XOR2_X1 _5899_ (.A(_1700_),
    .B(_1702_),
    .Z(_1703_));
 AND2_X1 _5900_ (.A1(_1699_),
    .A2(_1703_),
    .ZN(_1704_));
 AND2_X1 _5901_ (.A1(_1700_),
    .A2(_1702_),
    .ZN(_1705_));
 OAI21_X1 _5902_ (.A(_1698_),
    .B1(_1704_),
    .B2(_1705_),
    .ZN(_1706_));
 NAND2_X1 _5903_ (.A1(\fir.p6[9] ),
    .A2(\fir.p6[10] ),
    .ZN(_1707_));
 NAND2_X1 _5904_ (.A1(\fir.p7[8] ),
    .A2(\fir.p7[6] ),
    .ZN(_1708_));
 XOR2_X1 _5905_ (.A(\fir.p6[11] ),
    .B(\fir.p6[10] ),
    .Z(_1709_));
 XNOR2_X1 _5906_ (.A(_1708_),
    .B(_1709_),
    .ZN(_1710_));
 XOR2_X1 _5907_ (.A(_1707_),
    .B(_1710_),
    .Z(_1711_));
 NOR3_X1 _5908_ (.A1(_1705_),
    .A2(_1704_),
    .A3(_1698_),
    .ZN(_1712_));
 OAI21_X1 _5909_ (.A(_1706_),
    .B1(_1711_),
    .B2(_1712_),
    .ZN(_1713_));
 XOR2_X1 _5910_ (.A(_1662_),
    .B(_1674_),
    .Z(_1714_));
 NAND2_X1 _5911_ (.A1(_1713_),
    .A2(_1714_),
    .ZN(_1715_));
 NAND3_X1 _5912_ (.A1(\fir.p7[8] ),
    .A2(\fir.p7[6] ),
    .A3(_1709_),
    .ZN(_1716_));
 NAND3_X1 _5913_ (.A1(\fir.p6[9] ),
    .A2(\fir.p6[10] ),
    .A3(_1710_),
    .ZN(_1717_));
 NAND2_X1 _5914_ (.A1(_1716_),
    .A2(_1717_),
    .ZN(_1718_));
 XOR2_X1 _5915_ (.A(\fir.p6[6] ),
    .B(_1718_),
    .Z(_1719_));
 XOR2_X1 _5916_ (.A(_1713_),
    .B(_1714_),
    .Z(_1720_));
 NAND2_X1 _5917_ (.A1(_1719_),
    .A2(_1720_),
    .ZN(_1721_));
 NAND2_X1 _5918_ (.A1(_1715_),
    .A2(_1721_),
    .ZN(_1722_));
 XOR2_X1 _5919_ (.A(_1659_),
    .B(_1680_),
    .Z(_1723_));
 NAND2_X1 _5920_ (.A1(_1722_),
    .A2(_1723_),
    .ZN(_1724_));
 AND2_X1 _5921_ (.A1(\fir.p6[6] ),
    .A2(_1718_),
    .ZN(_1725_));
 XOR2_X1 _5922_ (.A(_1722_),
    .B(_1723_),
    .Z(_1726_));
 NAND2_X1 _5923_ (.A1(_1725_),
    .A2(_1726_),
    .ZN(_1727_));
 NAND2_X1 _5924_ (.A1(_1724_),
    .A2(_1727_),
    .ZN(_1728_));
 XOR2_X1 _5925_ (.A(_1686_),
    .B(_1687_),
    .Z(_1729_));
 AND2_X1 _5926_ (.A1(_1728_),
    .A2(_1729_),
    .ZN(_1730_));
 XOR2_X1 _5927_ (.A(_1689_),
    .B(_1690_),
    .Z(_1731_));
 NAND2_X1 _5928_ (.A1(_1730_),
    .A2(_1731_),
    .ZN(_1732_));
 XNOR2_X1 _5929_ (.A(_1730_),
    .B(_1731_),
    .ZN(_1733_));
 XOR2_X1 _5930_ (.A(\fir.p6[9] ),
    .B(\fir.p6[10] ),
    .Z(_1734_));
 NAND3_X1 _5931_ (.A1(\fir.p7[7] ),
    .A2(\fir.p7[5] ),
    .A3(_1734_),
    .ZN(_1735_));
 NAND2_X1 _5932_ (.A1(\fir.p7[7] ),
    .A2(\fir.p7[5] ),
    .ZN(_1736_));
 XNOR2_X1 _5933_ (.A(_1736_),
    .B(_1734_),
    .ZN(_1737_));
 NAND3_X1 _5934_ (.A1(\fir.p6[9] ),
    .A2(\fir.p6[8] ),
    .A3(_1737_),
    .ZN(_1738_));
 NAND2_X1 _5935_ (.A1(_1735_),
    .A2(_1738_),
    .ZN(_1739_));
 XOR2_X1 _5936_ (.A(_1699_),
    .B(_1703_),
    .Z(_1740_));
 XOR2_X1 _5937_ (.A(\fir.p7[7] ),
    .B(\fir.p7[5] ),
    .Z(_1741_));
 XNOR2_X1 _5938_ (.A(\fir.p7[9] ),
    .B(_1701_),
    .ZN(_1742_));
 XOR2_X1 _5939_ (.A(_0786_),
    .B(_0787_),
    .Z(_1743_));
 XNOR2_X1 _5940_ (.A(_1743_),
    .B(_0829_),
    .ZN(_1744_));
 NAND2_X1 _5941_ (.A1(\fir.p7[8] ),
    .A2(_1744_),
    .ZN(_1745_));
 XOR2_X1 _5942_ (.A(_1742_),
    .B(_1745_),
    .Z(_1746_));
 AND2_X1 _5943_ (.A1(_1741_),
    .A2(_1746_),
    .ZN(_1747_));
 NOR2_X1 _5944_ (.A1(_1742_),
    .A2(_1745_),
    .ZN(_1748_));
 OAI21_X1 _5945_ (.A(_1740_),
    .B1(_1747_),
    .B2(_1748_),
    .ZN(_1749_));
 NAND2_X1 _5946_ (.A1(\fir.p6[9] ),
    .A2(\fir.p6[8] ),
    .ZN(_1750_));
 XNOR2_X1 _5947_ (.A(_1750_),
    .B(_1737_),
    .ZN(_1751_));
 NOR2_X1 _5948_ (.A1(_1748_),
    .A2(_1747_),
    .ZN(_1752_));
 XNOR2_X1 _5949_ (.A(_1752_),
    .B(_1740_),
    .ZN(_1753_));
 NAND2_X1 _5950_ (.A1(_1751_),
    .A2(_1753_),
    .ZN(_1754_));
 NAND2_X1 _5951_ (.A1(_1749_),
    .A2(_1754_),
    .ZN(_1755_));
 NOR2_X1 _5952_ (.A1(_1705_),
    .A2(_1704_),
    .ZN(_1756_));
 XNOR2_X1 _5953_ (.A(_1756_),
    .B(_1698_),
    .ZN(_1757_));
 XNOR2_X1 _5954_ (.A(_1711_),
    .B(_1757_),
    .ZN(_1758_));
 AND2_X1 _5955_ (.A1(_1755_),
    .A2(_1758_),
    .ZN(_1759_));
 XOR2_X1 _5956_ (.A(\fir.p6[5] ),
    .B(_1739_),
    .Z(_1760_));
 XOR2_X1 _5957_ (.A(_1755_),
    .B(_1758_),
    .Z(_1761_));
 AOI21_X1 _5958_ (.A(_1759_),
    .B1(_1760_),
    .B2(_1761_),
    .ZN(_1762_));
 XNOR2_X1 _5959_ (.A(_1719_),
    .B(_1720_),
    .ZN(_1763_));
 XOR2_X1 _5960_ (.A(_1762_),
    .B(_1763_),
    .Z(_1764_));
 NAND3_X1 _5961_ (.A1(\fir.p6[5] ),
    .A2(_1739_),
    .A3(_1764_),
    .ZN(_1765_));
 OAI21_X1 _5962_ (.A(_1765_),
    .B1(_1763_),
    .B2(_1762_),
    .ZN(_1766_));
 XOR2_X1 _5963_ (.A(_1725_),
    .B(_1726_),
    .Z(_1767_));
 XOR2_X1 _5964_ (.A(_1728_),
    .B(_1729_),
    .Z(_1768_));
 AND3_X1 _5965_ (.A1(_1766_),
    .A2(_1767_),
    .A3(_1768_),
    .ZN(_1769_));
 NAND2_X1 _5966_ (.A1(_1766_),
    .A2(_1767_),
    .ZN(_1770_));
 XNOR2_X1 _5967_ (.A(_1770_),
    .B(_1768_),
    .ZN(_1771_));
 XOR2_X1 _5968_ (.A(\fir.p7[8] ),
    .B(_1744_),
    .Z(_1772_));
 XOR2_X1 _5969_ (.A(_0824_),
    .B(_0827_),
    .Z(_1773_));
 AND2_X1 _5970_ (.A1(\fir.p7[7] ),
    .A2(_1773_),
    .ZN(_1774_));
 NAND2_X1 _5971_ (.A1(_1772_),
    .A2(_1774_),
    .ZN(_1775_));
 XOR2_X1 _5972_ (.A(\fir.p7[6] ),
    .B(\fir.p7[4] ),
    .Z(_1776_));
 XOR2_X1 _5973_ (.A(_1772_),
    .B(_1774_),
    .Z(_1777_));
 NAND2_X1 _5974_ (.A1(_1776_),
    .A2(_1777_),
    .ZN(_1778_));
 NAND2_X1 _5975_ (.A1(_1775_),
    .A2(_1778_),
    .ZN(_1779_));
 XOR2_X1 _5976_ (.A(_1741_),
    .B(_1746_),
    .Z(_1780_));
 NAND2_X1 _5977_ (.A1(_1779_),
    .A2(_1780_),
    .ZN(_1781_));
 NAND2_X1 _5978_ (.A1(\fir.p6[8] ),
    .A2(\fir.p6[7] ),
    .ZN(_1782_));
 NAND2_X1 _5979_ (.A1(\fir.p7[6] ),
    .A2(\fir.p7[4] ),
    .ZN(_1783_));
 XOR2_X1 _5980_ (.A(\fir.p6[9] ),
    .B(\fir.p6[8] ),
    .Z(_1784_));
 XNOR2_X1 _5981_ (.A(_1783_),
    .B(_1784_),
    .ZN(_1785_));
 XNOR2_X1 _5982_ (.A(_1782_),
    .B(_1785_),
    .ZN(_1786_));
 XOR2_X1 _5983_ (.A(_1779_),
    .B(_1780_),
    .Z(_1787_));
 NAND2_X1 _5984_ (.A1(_1786_),
    .A2(_1787_),
    .ZN(_1788_));
 NAND2_X1 _5985_ (.A1(_1781_),
    .A2(_1788_),
    .ZN(_1789_));
 XOR2_X1 _5986_ (.A(_1751_),
    .B(_1753_),
    .Z(_1790_));
 NAND2_X1 _5987_ (.A1(_1789_),
    .A2(_1790_),
    .ZN(_1791_));
 NAND3_X1 _5988_ (.A1(\fir.p7[6] ),
    .A2(\fir.p7[4] ),
    .A3(_1784_),
    .ZN(_1792_));
 NAND3_X1 _5989_ (.A1(\fir.p6[8] ),
    .A2(\fir.p6[7] ),
    .A3(_1785_),
    .ZN(_1793_));
 NAND2_X1 _5990_ (.A1(_1792_),
    .A2(_1793_),
    .ZN(_1794_));
 XOR2_X1 _5991_ (.A(\fir.p6[4] ),
    .B(_1794_),
    .Z(_1795_));
 XOR2_X1 _5992_ (.A(_1789_),
    .B(_1790_),
    .Z(_1796_));
 NAND2_X1 _5993_ (.A1(_1795_),
    .A2(_1796_),
    .ZN(_1797_));
 NAND2_X1 _5994_ (.A1(_1791_),
    .A2(_1797_),
    .ZN(_1798_));
 XOR2_X1 _5995_ (.A(_1760_),
    .B(_1761_),
    .Z(_1799_));
 NAND2_X1 _5996_ (.A1(_1798_),
    .A2(_1799_),
    .ZN(_1800_));
 AND2_X1 _5997_ (.A1(\fir.p6[4] ),
    .A2(_1794_),
    .ZN(_1801_));
 XOR2_X1 _5998_ (.A(_1798_),
    .B(_1799_),
    .Z(_1802_));
 NAND2_X1 _5999_ (.A1(_1801_),
    .A2(_1802_),
    .ZN(_1803_));
 NAND2_X1 _6000_ (.A1(_1800_),
    .A2(_1803_),
    .ZN(_1804_));
 NAND2_X1 _6001_ (.A1(\fir.p6[5] ),
    .A2(_1739_),
    .ZN(_1805_));
 XNOR2_X1 _6002_ (.A(_1805_),
    .B(_1764_),
    .ZN(_1806_));
 XOR2_X1 _6003_ (.A(_1766_),
    .B(_1767_),
    .Z(_1807_));
 NAND3_X1 _6004_ (.A1(_1804_),
    .A2(_1806_),
    .A3(_1807_),
    .ZN(_1808_));
 NAND2_X1 _6005_ (.A1(_1804_),
    .A2(_1806_),
    .ZN(_1809_));
 XNOR2_X1 _6006_ (.A(_1809_),
    .B(_1807_),
    .ZN(_1810_));
 INV_X1 _6007_ (.A(_1810_),
    .ZN(_1811_));
 XOR2_X1 _6008_ (.A(_1804_),
    .B(_1806_),
    .Z(_1812_));
 XOR2_X1 _6009_ (.A(\fir.p6[8] ),
    .B(\fir.p6[7] ),
    .Z(_1813_));
 NAND3_X1 _6010_ (.A1(\fir.p7[3] ),
    .A2(\fir.p7[5] ),
    .A3(_1813_),
    .ZN(_1814_));
 NAND2_X1 _6011_ (.A1(\fir.p7[3] ),
    .A2(\fir.p7[5] ),
    .ZN(_1815_));
 XNOR2_X1 _6012_ (.A(_1815_),
    .B(_1813_),
    .ZN(_1816_));
 NAND3_X1 _6013_ (.A1(\fir.p6[7] ),
    .A2(\fir.p6[6] ),
    .A3(_1816_),
    .ZN(_1817_));
 NAND2_X1 _6014_ (.A1(_1814_),
    .A2(_1817_),
    .ZN(_1818_));
 XOR2_X1 _6015_ (.A(\fir.p7[3] ),
    .B(\fir.p7[5] ),
    .Z(_1819_));
 XNOR2_X1 _6016_ (.A(\fir.p7[7] ),
    .B(_1773_),
    .ZN(_1820_));
 INV_X1 _6017_ (.A(\fir.p7[6] ),
    .ZN(_1821_));
 XNOR2_X1 _6018_ (.A(_0820_),
    .B(_0823_),
    .ZN(_1822_));
 NOR2_X1 _6019_ (.A1(_1821_),
    .A2(_1822_),
    .ZN(_1823_));
 XNOR2_X1 _6020_ (.A(_1820_),
    .B(_1823_),
    .ZN(_1824_));
 NAND2_X1 _6021_ (.A1(_1819_),
    .A2(_1824_),
    .ZN(_1825_));
 INV_X1 _6022_ (.A(_1823_),
    .ZN(_1826_));
 OAI21_X1 _6023_ (.A(_1825_),
    .B1(_1826_),
    .B2(_1820_),
    .ZN(_1827_));
 XOR2_X1 _6024_ (.A(_1776_),
    .B(_1777_),
    .Z(_1828_));
 NAND2_X1 _6025_ (.A1(_1827_),
    .A2(_1828_),
    .ZN(_1829_));
 NAND2_X1 _6026_ (.A1(\fir.p6[7] ),
    .A2(\fir.p6[6] ),
    .ZN(_1830_));
 XNOR2_X1 _6027_ (.A(_1830_),
    .B(_1816_),
    .ZN(_1831_));
 XOR2_X1 _6028_ (.A(_1827_),
    .B(_1828_),
    .Z(_1832_));
 NAND2_X1 _6029_ (.A1(_1831_),
    .A2(_1832_),
    .ZN(_1833_));
 NAND2_X1 _6030_ (.A1(_1829_),
    .A2(_1833_),
    .ZN(_1834_));
 XOR2_X1 _6031_ (.A(_1786_),
    .B(_1787_),
    .Z(_1835_));
 AND2_X1 _6032_ (.A1(_1834_),
    .A2(_1835_),
    .ZN(_1836_));
 XOR2_X1 _6033_ (.A(\fir.p6[3] ),
    .B(_1818_),
    .Z(_1837_));
 XOR2_X1 _6034_ (.A(_1834_),
    .B(_1835_),
    .Z(_1838_));
 AOI21_X1 _6035_ (.A(_1836_),
    .B1(_1837_),
    .B2(_1838_),
    .ZN(_1839_));
 XNOR2_X1 _6036_ (.A(_1795_),
    .B(_1796_),
    .ZN(_1840_));
 XOR2_X1 _6037_ (.A(_1839_),
    .B(_1840_),
    .Z(_1841_));
 NAND3_X1 _6038_ (.A1(\fir.p6[3] ),
    .A2(_1818_),
    .A3(_1841_),
    .ZN(_1842_));
 OAI21_X1 _6039_ (.A(_1842_),
    .B1(_1840_),
    .B2(_1839_),
    .ZN(_1843_));
 XOR2_X1 _6040_ (.A(_1801_),
    .B(_1802_),
    .Z(_1844_));
 AND2_X1 _6041_ (.A1(_1843_),
    .A2(_1844_),
    .ZN(_1845_));
 AND2_X1 _6042_ (.A1(_1812_),
    .A2(_1845_),
    .ZN(_1846_));
 XOR2_X1 _6043_ (.A(_1812_),
    .B(_1845_),
    .Z(_1847_));
 XOR2_X1 _6044_ (.A(\fir.p7[2] ),
    .B(\fir.p7[4] ),
    .Z(_1848_));
 XNOR2_X1 _6045_ (.A(_1821_),
    .B(_1822_),
    .ZN(_1849_));
 XOR2_X1 _6046_ (.A(_0817_),
    .B(_0818_),
    .Z(_1850_));
 NAND2_X1 _6047_ (.A1(\fir.p7[5] ),
    .A2(_1850_),
    .ZN(_1851_));
 XOR2_X1 _6048_ (.A(_1849_),
    .B(_1851_),
    .Z(_1852_));
 NAND2_X1 _6049_ (.A1(_1848_),
    .A2(_1852_),
    .ZN(_1853_));
 OAI21_X1 _6050_ (.A(_1853_),
    .B1(_1851_),
    .B2(_1849_),
    .ZN(_1854_));
 XOR2_X1 _6051_ (.A(_1819_),
    .B(_1824_),
    .Z(_1855_));
 NAND2_X1 _6052_ (.A1(_1854_),
    .A2(_1855_),
    .ZN(_1856_));
 NAND2_X1 _6053_ (.A1(\fir.p6[6] ),
    .A2(\fir.p6[5] ),
    .ZN(_1857_));
 NAND2_X1 _6054_ (.A1(\fir.p7[2] ),
    .A2(\fir.p7[4] ),
    .ZN(_1858_));
 XOR2_X1 _6055_ (.A(\fir.p6[7] ),
    .B(\fir.p6[6] ),
    .Z(_1859_));
 XNOR2_X1 _6056_ (.A(_1858_),
    .B(_1859_),
    .ZN(_1860_));
 XNOR2_X1 _6057_ (.A(_1857_),
    .B(_1860_),
    .ZN(_1861_));
 XOR2_X1 _6058_ (.A(_1854_),
    .B(_1855_),
    .Z(_1862_));
 NAND2_X1 _6059_ (.A1(_1861_),
    .A2(_1862_),
    .ZN(_1863_));
 NAND2_X1 _6060_ (.A1(_1856_),
    .A2(_1863_),
    .ZN(_1864_));
 XOR2_X1 _6061_ (.A(_1831_),
    .B(_1832_),
    .Z(_1865_));
 NAND2_X1 _6062_ (.A1(_1864_),
    .A2(_1865_),
    .ZN(_1866_));
 NAND3_X1 _6063_ (.A1(\fir.p7[2] ),
    .A2(\fir.p7[4] ),
    .A3(_1859_),
    .ZN(_1867_));
 NAND3_X1 _6064_ (.A1(\fir.p6[6] ),
    .A2(\fir.p6[5] ),
    .A3(_1860_),
    .ZN(_1868_));
 NAND2_X1 _6065_ (.A1(_1867_),
    .A2(_1868_),
    .ZN(_1869_));
 XOR2_X1 _6066_ (.A(\fir.p6[2] ),
    .B(_1869_),
    .Z(_1870_));
 XOR2_X1 _6067_ (.A(_1864_),
    .B(_1865_),
    .Z(_1871_));
 NAND2_X1 _6068_ (.A1(_1870_),
    .A2(_1871_),
    .ZN(_1872_));
 NAND2_X1 _6069_ (.A1(_1866_),
    .A2(_1872_),
    .ZN(_1873_));
 XOR2_X1 _6070_ (.A(_1837_),
    .B(_1838_),
    .Z(_1874_));
 NAND2_X1 _6071_ (.A1(_1873_),
    .A2(_1874_),
    .ZN(_1875_));
 AND2_X1 _6072_ (.A1(\fir.p6[2] ),
    .A2(_1869_),
    .ZN(_1876_));
 XOR2_X1 _6073_ (.A(_1873_),
    .B(_1874_),
    .Z(_1877_));
 NAND2_X1 _6074_ (.A1(_1876_),
    .A2(_1877_),
    .ZN(_1878_));
 NAND2_X1 _6075_ (.A1(_1875_),
    .A2(_1878_),
    .ZN(_1879_));
 NAND2_X1 _6076_ (.A1(\fir.p6[3] ),
    .A2(_1818_),
    .ZN(_1880_));
 XNOR2_X1 _6077_ (.A(_1880_),
    .B(_1841_),
    .ZN(_1881_));
 AND2_X1 _6078_ (.A1(_1879_),
    .A2(_1881_),
    .ZN(_1882_));
 XOR2_X1 _6079_ (.A(_1843_),
    .B(_1844_),
    .Z(_1883_));
 NAND2_X1 _6080_ (.A1(_1882_),
    .A2(_1883_),
    .ZN(_1884_));
 XNOR2_X1 _6081_ (.A(_1882_),
    .B(_1883_),
    .ZN(_1885_));
 NAND2_X1 _6082_ (.A1(\fir.p6[5] ),
    .A2(\fir.p6[4] ),
    .ZN(_1886_));
 NAND2_X1 _6083_ (.A1(\fir.p7[1] ),
    .A2(\fir.p7[3] ),
    .ZN(_1887_));
 XOR2_X1 _6084_ (.A(\fir.p6[6] ),
    .B(\fir.p6[5] ),
    .Z(_1888_));
 XNOR2_X1 _6085_ (.A(_1887_),
    .B(_1888_),
    .ZN(_1889_));
 XNOR2_X1 _6086_ (.A(_1886_),
    .B(_1889_),
    .ZN(_1890_));
 XNOR2_X1 _6087_ (.A(\fir.p7[5] ),
    .B(_1850_),
    .ZN(_1891_));
 XOR2_X1 _6088_ (.A(_0814_),
    .B(_0816_),
    .Z(_1892_));
 NAND2_X1 _6089_ (.A1(\fir.p7[4] ),
    .A2(_1892_),
    .ZN(_1893_));
 NOR2_X1 _6090_ (.A1(_1891_),
    .A2(_1893_),
    .ZN(_1894_));
 XOR2_X1 _6091_ (.A(\fir.p7[1] ),
    .B(\fir.p7[3] ),
    .Z(_1895_));
 XOR2_X1 _6092_ (.A(_1891_),
    .B(_1893_),
    .Z(_1896_));
 AOI21_X1 _6093_ (.A(_1894_),
    .B1(_1895_),
    .B2(_1896_),
    .ZN(_1897_));
 XNOR2_X1 _6094_ (.A(_1848_),
    .B(_1852_),
    .ZN(_1898_));
 XOR2_X1 _6095_ (.A(_1897_),
    .B(_1898_),
    .Z(_1899_));
 NAND2_X1 _6096_ (.A1(_1890_),
    .A2(_1899_),
    .ZN(_1900_));
 OAI21_X1 _6097_ (.A(_1900_),
    .B1(_1898_),
    .B2(_1897_),
    .ZN(_1901_));
 XOR2_X1 _6098_ (.A(_1861_),
    .B(_1862_),
    .Z(_1902_));
 NAND2_X1 _6099_ (.A1(_1901_),
    .A2(_1902_),
    .ZN(_1903_));
 INV_X1 _6100_ (.A(net213),
    .ZN(_1904_));
 NAND3_X1 _6101_ (.A1(\fir.p7[1] ),
    .A2(\fir.p7[3] ),
    .A3(_1888_),
    .ZN(_1905_));
 NAND3_X1 _6102_ (.A1(\fir.p6[5] ),
    .A2(\fir.p6[4] ),
    .A3(_1889_),
    .ZN(_1906_));
 NAND2_X1 _6103_ (.A1(_1905_),
    .A2(_1906_),
    .ZN(_1907_));
 XNOR2_X1 _6104_ (.A(_1904_),
    .B(_1907_),
    .ZN(_1908_));
 XOR2_X1 _6105_ (.A(_1901_),
    .B(_1902_),
    .Z(_1909_));
 NAND2_X1 _6106_ (.A1(_1908_),
    .A2(_1909_),
    .ZN(_1910_));
 NAND2_X1 _6107_ (.A1(_1903_),
    .A2(_1910_),
    .ZN(_1911_));
 XOR2_X1 _6108_ (.A(_1870_),
    .B(_1871_),
    .Z(_1912_));
 NAND2_X1 _6109_ (.A1(_1911_),
    .A2(_1912_),
    .ZN(_1913_));
 AOI21_X1 _6110_ (.A(_1904_),
    .B1(_1905_),
    .B2(_1906_),
    .ZN(_1914_));
 XOR2_X1 _6111_ (.A(_1911_),
    .B(_1912_),
    .Z(_1915_));
 NAND2_X1 _6112_ (.A1(_1914_),
    .A2(_1915_),
    .ZN(_1916_));
 NAND2_X1 _6113_ (.A1(_1913_),
    .A2(_1916_),
    .ZN(_1917_));
 XOR2_X1 _6114_ (.A(_1876_),
    .B(_1877_),
    .Z(_1918_));
 AND2_X1 _6115_ (.A1(_1917_),
    .A2(_1918_),
    .ZN(_1919_));
 XOR2_X1 _6116_ (.A(_1879_),
    .B(_1881_),
    .Z(_1920_));
 AND2_X1 _6117_ (.A1(_1919_),
    .A2(_1920_),
    .ZN(_1921_));
 XOR2_X1 _6118_ (.A(_1919_),
    .B(_1920_),
    .Z(_1922_));
 XNOR2_X1 _6119_ (.A(_1914_),
    .B(_1915_),
    .ZN(_1923_));
 INV_X1 _6120_ (.A(net120),
    .ZN(_1924_));
 XOR2_X1 _6121_ (.A(\fir.p6[5] ),
    .B(\fir.p6[4] ),
    .Z(_1925_));
 NAND3_X1 _6122_ (.A1(\fir.p7[0] ),
    .A2(\fir.p7[2] ),
    .A3(_1925_),
    .ZN(_1926_));
 NAND2_X1 _6123_ (.A1(\fir.p7[0] ),
    .A2(\fir.p7[2] ),
    .ZN(_1927_));
 XNOR2_X1 _6124_ (.A(_1927_),
    .B(_1925_),
    .ZN(_1928_));
 NAND3_X1 _6125_ (.A1(\fir.p6[4] ),
    .A2(\fir.p6[3] ),
    .A3(_1928_),
    .ZN(_1929_));
 AOI21_X1 _6126_ (.A(_1924_),
    .B1(_1926_),
    .B2(_1929_),
    .ZN(_1930_));
 XOR2_X1 _6127_ (.A(\fir.p7[0] ),
    .B(\fir.p7[2] ),
    .Z(_1931_));
 XNOR2_X1 _6128_ (.A(\fir.p7[4] ),
    .B(_1892_),
    .ZN(_1932_));
 NOR2_X1 _6129_ (.A1(_0811_),
    .A2(_0812_),
    .ZN(_1933_));
 XNOR2_X1 _6130_ (.A(_1933_),
    .B(_0813_),
    .ZN(_1934_));
 NAND2_X1 _6131_ (.A1(\fir.p7[3] ),
    .A2(_1934_),
    .ZN(_1935_));
 XOR2_X1 _6132_ (.A(_1932_),
    .B(_1935_),
    .Z(_1936_));
 NAND2_X1 _6133_ (.A1(_1931_),
    .A2(_1936_),
    .ZN(_1937_));
 OAI21_X1 _6134_ (.A(_1937_),
    .B1(_1935_),
    .B2(_1932_),
    .ZN(_1938_));
 XOR2_X1 _6135_ (.A(_1895_),
    .B(_1896_),
    .Z(_1939_));
 NAND2_X1 _6136_ (.A1(\fir.p6[4] ),
    .A2(\fir.p6[3] ),
    .ZN(_1940_));
 XNOR2_X1 _6137_ (.A(_1940_),
    .B(_1928_),
    .ZN(_1941_));
 XOR2_X1 _6138_ (.A(_1938_),
    .B(_1939_),
    .Z(_1942_));
 AOI22_X1 _6139_ (.A1(_1938_),
    .A2(_1939_),
    .B1(_1941_),
    .B2(_1942_),
    .ZN(_1943_));
 XNOR2_X1 _6140_ (.A(_1890_),
    .B(_1899_),
    .ZN(_1944_));
 NOR2_X1 _6141_ (.A1(_1943_),
    .A2(_1944_),
    .ZN(_1945_));
 NAND2_X1 _6142_ (.A1(_1926_),
    .A2(_1929_),
    .ZN(_1946_));
 XNOR2_X1 _6143_ (.A(\fir.p6[0] ),
    .B(_1946_),
    .ZN(_1947_));
 XNOR2_X1 _6144_ (.A(_1943_),
    .B(_1944_),
    .ZN(_1948_));
 NOR2_X1 _6145_ (.A1(_1947_),
    .A2(_1948_),
    .ZN(_1949_));
 NOR2_X1 _6146_ (.A1(_1945_),
    .A2(_1949_),
    .ZN(_1950_));
 XOR2_X1 _6147_ (.A(_1908_),
    .B(_1909_),
    .Z(_1951_));
 XNOR2_X1 _6148_ (.A(_1950_),
    .B(_1951_),
    .ZN(_1952_));
 NAND2_X1 _6149_ (.A1(_1930_),
    .A2(_1952_),
    .ZN(_1953_));
 OAI21_X1 _6150_ (.A(_1951_),
    .B1(_1949_),
    .B2(_1945_),
    .ZN(_1954_));
 AOI21_X1 _6151_ (.A(_1923_),
    .B1(_1953_),
    .B2(_1954_),
    .ZN(_1955_));
 XOR2_X1 _6152_ (.A(_1917_),
    .B(_1918_),
    .Z(_1956_));
 NAND2_X1 _6153_ (.A1(_1955_),
    .A2(_1956_),
    .ZN(_1957_));
 XNOR2_X1 _6154_ (.A(_1955_),
    .B(_1956_),
    .ZN(_1958_));
 NAND3_X1 _6155_ (.A1(_1954_),
    .A2(_1953_),
    .A3(_1923_),
    .ZN(_1959_));
 AND2_X1 _6156_ (.A1(_1947_),
    .A2(_1948_),
    .ZN(_1960_));
 XNOR2_X1 _6157_ (.A(_1941_),
    .B(_1942_),
    .ZN(_1961_));
 NAND2_X1 _6158_ (.A1(\fir.p6[3] ),
    .A2(\fir.p6[2] ),
    .ZN(_1962_));
 XOR2_X1 _6159_ (.A(\fir.p6[4] ),
    .B(\fir.p6[3] ),
    .Z(_1963_));
 XNOR2_X1 _6160_ (.A(_1962_),
    .B(_1963_),
    .ZN(_1964_));
 XOR2_X1 _6161_ (.A(_1931_),
    .B(_1936_),
    .Z(_1965_));
 XNOR2_X1 _6162_ (.A(\fir.p7[3] ),
    .B(_1934_),
    .ZN(_1966_));
 XOR2_X1 _6163_ (.A(_0811_),
    .B(_0812_),
    .Z(_1967_));
 NAND2_X1 _6164_ (.A1(\fir.p7[2] ),
    .A2(_1967_),
    .ZN(_1968_));
 XOR2_X1 _6165_ (.A(_1966_),
    .B(_1968_),
    .Z(_1969_));
 AND2_X1 _6166_ (.A1(\fir.p7[1] ),
    .A2(_1969_),
    .ZN(_1970_));
 NOR2_X1 _6167_ (.A1(_1966_),
    .A2(_1968_),
    .ZN(_1971_));
 OAI21_X1 _6168_ (.A(_1965_),
    .B1(_1970_),
    .B2(_1971_),
    .ZN(_1972_));
 OR3_X1 _6169_ (.A1(_1971_),
    .A2(_1970_),
    .A3(_1965_),
    .ZN(_1973_));
 AND2_X1 _6170_ (.A1(_1972_),
    .A2(_1973_),
    .ZN(_1974_));
 NAND2_X1 _6171_ (.A1(_1964_),
    .A2(_1974_),
    .ZN(_1975_));
 AOI21_X1 _6172_ (.A(_1961_),
    .B1(_1975_),
    .B2(_1972_),
    .ZN(_1976_));
 NOR2_X1 _6173_ (.A1(\fir.p6[4] ),
    .A2(_1962_),
    .ZN(_1977_));
 AND3_X1 _6174_ (.A1(_1972_),
    .A2(_1975_),
    .A3(_1961_),
    .ZN(_1978_));
 NOR2_X1 _6175_ (.A1(_1976_),
    .A2(_1978_),
    .ZN(_1979_));
 XOR2_X1 _6176_ (.A(_1977_),
    .B(_1979_),
    .Z(_1980_));
 NAND2_X1 _6177_ (.A1(\fir.p6[2] ),
    .A2(\fir.p6[1] ),
    .ZN(_1981_));
 NOR2_X1 _6178_ (.A1(\fir.p6[3] ),
    .A2(_1981_),
    .ZN(_1982_));
 XNOR2_X1 _6179_ (.A(\fir.p7[1] ),
    .B(_1969_),
    .ZN(_1983_));
 XNOR2_X1 _6180_ (.A(\fir.p7[2] ),
    .B(_1967_),
    .ZN(_1984_));
 XNOR2_X1 _6181_ (.A(\fir.p5[0] ),
    .B(_0810_),
    .ZN(_1985_));
 INV_X1 _6182_ (.A(_1985_),
    .ZN(_1986_));
 NAND2_X1 _6183_ (.A1(\fir.p7[1] ),
    .A2(_1986_),
    .ZN(_1987_));
 XOR2_X1 _6184_ (.A(_1984_),
    .B(_1987_),
    .Z(_1988_));
 NAND2_X1 _6185_ (.A1(\fir.p7[0] ),
    .A2(_1988_),
    .ZN(_1989_));
 OR2_X1 _6186_ (.A1(_1984_),
    .A2(_1987_),
    .ZN(_1990_));
 AOI21_X1 _6187_ (.A(_1983_),
    .B1(_1989_),
    .B2(_1990_),
    .ZN(_1991_));
 XOR2_X1 _6188_ (.A(\fir.p6[3] ),
    .B(\fir.p6[2] ),
    .Z(_1992_));
 XNOR2_X1 _6189_ (.A(_1981_),
    .B(_1992_),
    .ZN(_1993_));
 AND3_X1 _6190_ (.A1(_1990_),
    .A2(_1989_),
    .A3(_1983_),
    .ZN(_1994_));
 NOR2_X1 _6191_ (.A1(_1991_),
    .A2(_1994_),
    .ZN(_1995_));
 AOI21_X1 _6192_ (.A(_1991_),
    .B1(_1993_),
    .B2(_1995_),
    .ZN(_1996_));
 XNOR2_X1 _6193_ (.A(_1964_),
    .B(_1974_),
    .ZN(_1997_));
 XOR2_X1 _6194_ (.A(_1996_),
    .B(_1997_),
    .Z(_1998_));
 NAND2_X1 _6195_ (.A1(_1982_),
    .A2(_1998_),
    .ZN(_1999_));
 NOR2_X1 _6196_ (.A1(_1982_),
    .A2(_1998_),
    .ZN(_2000_));
 XOR2_X1 _6197_ (.A(_1993_),
    .B(_1995_),
    .Z(_2001_));
 NAND2_X1 _6198_ (.A1(\fir.p6[1] ),
    .A2(\fir.p6[0] ),
    .ZN(_2002_));
 XNOR2_X1 _6199_ (.A(\fir.p6[2] ),
    .B(\fir.p6[1] ),
    .ZN(_2003_));
 XNOR2_X1 _6200_ (.A(_2002_),
    .B(_2003_),
    .ZN(_2004_));
 XNOR2_X1 _6201_ (.A(\fir.p3[0] ),
    .B(_3490_),
    .ZN(_2005_));
 NAND2_X1 _6202_ (.A1(\fir.p7[0] ),
    .A2(_2005_),
    .ZN(_2006_));
 XOR2_X1 _6203_ (.A(\fir.p7[1] ),
    .B(_1985_),
    .Z(_2007_));
 NOR2_X1 _6204_ (.A1(_2006_),
    .A2(_2007_),
    .ZN(_2008_));
 XNOR2_X1 _6205_ (.A(\fir.p7[0] ),
    .B(_1988_),
    .ZN(_2009_));
 XOR2_X1 _6206_ (.A(_2008_),
    .B(_2009_),
    .Z(_2010_));
 NOR2_X1 _6207_ (.A1(_2004_),
    .A2(_2010_),
    .ZN(_2011_));
 NOR3_X1 _6208_ (.A1(_2006_),
    .A2(_2007_),
    .A3(_2009_),
    .ZN(_2012_));
 OAI21_X1 _6209_ (.A(_2001_),
    .B1(_2011_),
    .B2(_2012_),
    .ZN(_2013_));
 OR3_X1 _6210_ (.A1(_2012_),
    .A2(_2011_),
    .A3(_2001_),
    .ZN(_2014_));
 NAND2_X1 _6211_ (.A1(_2013_),
    .A2(_2014_),
    .ZN(_2015_));
 OR3_X1 _6212_ (.A1(\fir.p6[2] ),
    .A2(_2002_),
    .A3(_2015_),
    .ZN(_2016_));
 OAI211_X1 _6213_ (.A(_1904_),
    .B(\fir.p6[0] ),
    .C1(\fir.p7[0] ),
    .C2(_2005_),
    .ZN(_2017_));
 AND3_X1 _6214_ (.A1(_2006_),
    .A2(_2007_),
    .A3(_2017_),
    .ZN(_2018_));
 XNOR2_X1 _6215_ (.A(\fir.p7[0] ),
    .B(_2005_),
    .ZN(_2019_));
 NAND3_X1 _6216_ (.A1(\fir.p6[1] ),
    .A2(\fir.p6[0] ),
    .A3(_2019_),
    .ZN(_2020_));
 OAI221_X1 _6217_ (.A(_2020_),
    .B1(_2007_),
    .B2(_2006_),
    .C1(\fir.p6[1] ),
    .C2(\fir.p6[0] ),
    .ZN(_2021_));
 AOI211_X1 _6218_ (.A(_2018_),
    .B(_2021_),
    .C1(_2009_),
    .C2(_2004_),
    .ZN(_2022_));
 OAI21_X1 _6219_ (.A(_2015_),
    .B1(_2002_),
    .B2(\fir.p6[2] ),
    .ZN(_2023_));
 OAI211_X1 _6220_ (.A(_2022_),
    .B(_2023_),
    .C1(_2004_),
    .C2(_2010_),
    .ZN(_2024_));
 AND3_X1 _6221_ (.A1(_2013_),
    .A2(_2016_),
    .A3(_2024_),
    .ZN(_2025_));
 OAI221_X1 _6222_ (.A(_1999_),
    .B1(_2000_),
    .B2(_2025_),
    .C1(_1997_),
    .C2(_1996_),
    .ZN(_2026_));
 AOI221_X1 _6223_ (.A(_1976_),
    .B1(_1980_),
    .B2(_2026_),
    .C1(_1979_),
    .C2(_1977_),
    .ZN(_2027_));
 XNOR2_X1 _6224_ (.A(_1930_),
    .B(_1952_),
    .ZN(_2028_));
 NOR4_X1 _6225_ (.A1(_1949_),
    .A2(_1960_),
    .A3(_2027_),
    .A4(_2028_),
    .ZN(_2029_));
 NAND2_X1 _6226_ (.A1(_1959_),
    .A2(_2029_),
    .ZN(_2030_));
 OAI21_X1 _6227_ (.A(_1957_),
    .B1(_1958_),
    .B2(_2030_),
    .ZN(_2031_));
 AOI21_X1 _6228_ (.A(_1921_),
    .B1(_1922_),
    .B2(_2031_),
    .ZN(_2032_));
 OAI21_X1 _6229_ (.A(_1884_),
    .B1(_1885_),
    .B2(_2032_),
    .ZN(_2033_));
 AOI21_X1 _6230_ (.A(_1846_),
    .B1(_1847_),
    .B2(_2033_),
    .ZN(_2034_));
 OAI21_X1 _6231_ (.A(_1808_),
    .B1(_1811_),
    .B2(_2034_),
    .ZN(_2035_));
 AOI21_X1 _6232_ (.A(_1769_),
    .B1(_1771_),
    .B2(_2035_),
    .ZN(_2036_));
 OAI21_X1 _6233_ (.A(_1732_),
    .B1(_1733_),
    .B2(_2036_),
    .ZN(_2037_));
 AOI221_X1 _6234_ (.A(_1657_),
    .B1(_1694_),
    .B2(_1695_),
    .C1(_1697_),
    .C2(_2037_),
    .ZN(_2038_));
 XNOR2_X1 _6235_ (.A(_1628_),
    .B(_2038_),
    .ZN(_2039_));
 XOR2_X1 _6236_ (.A(_2037_),
    .B(_1696_),
    .Z(_2040_));
 XOR2_X1 _6237_ (.A(_1733_),
    .B(_2036_),
    .Z(_2041_));
 XOR2_X1 _6238_ (.A(_1771_),
    .B(_2035_),
    .Z(_2042_));
 XOR2_X1 _6239_ (.A(_1847_),
    .B(_2033_),
    .Z(_2043_));
 XOR2_X1 _6240_ (.A(_1958_),
    .B(_2030_),
    .Z(_2044_));
 XOR2_X1 _6241_ (.A(_1922_),
    .B(_2031_),
    .Z(_2045_));
 XOR2_X1 _6242_ (.A(_1885_),
    .B(_2032_),
    .Z(_2046_));
 AND3_X1 _6243_ (.A1(_2044_),
    .A2(_2045_),
    .A3(_2046_),
    .ZN(_2047_));
 NAND2_X1 _6244_ (.A1(_2043_),
    .A2(_2047_),
    .ZN(_2048_));
 XNOR2_X1 _6245_ (.A(_1811_),
    .B(_2034_),
    .ZN(_2049_));
 NOR2_X1 _6246_ (.A1(_2048_),
    .A2(_2049_),
    .ZN(_2050_));
 AND2_X1 _6247_ (.A1(_2042_),
    .A2(_2050_),
    .ZN(_2051_));
 AND2_X1 _6248_ (.A1(_2041_),
    .A2(_2051_),
    .ZN(_2052_));
 AND2_X1 _6249_ (.A1(_2040_),
    .A2(_2052_),
    .ZN(_2053_));
 AOI21_X1 _6250_ (.A(_1694_),
    .B1(_2037_),
    .B2(_1696_),
    .ZN(_2054_));
 XNOR2_X1 _6251_ (.A(_2054_),
    .B(_1695_),
    .ZN(_2055_));
 NAND3_X1 _6252_ (.A1(_2039_),
    .A2(_2053_),
    .A3(_2055_),
    .ZN(_2056_));
 NOR2_X1 _6253_ (.A1(_1535_),
    .A2(_1626_),
    .ZN(_2057_));
 AND2_X1 _6254_ (.A1(_1539_),
    .A2(_1624_),
    .ZN(_2058_));
 AOI21_X1 _6255_ (.A(_2058_),
    .B1(_1625_),
    .B2(_1537_),
    .ZN(_2059_));
 INV_X1 _6256_ (.A(_1621_),
    .ZN(_2060_));
 NOR2_X1 _6257_ (.A1(_1536_),
    .A2(\fir.p7[11] ),
    .ZN(_2061_));
 AOI21_X1 _6258_ (.A(_2060_),
    .B1(_1623_),
    .B2(_2061_),
    .ZN(_2062_));
 NOR2_X1 _6259_ (.A1(_1315_),
    .A2(_1617_),
    .ZN(_2063_));
 AND3_X1 _6260_ (.A1(_0991_),
    .A2(_1415_),
    .A3(_1523_),
    .ZN(_2064_));
 AOI21_X1 _6261_ (.A(_2063_),
    .B1(_1616_),
    .B2(_2064_),
    .ZN(_2065_));
 AND4_X1 _6262_ (.A1(_0991_),
    .A2(_1521_),
    .A3(_1522_),
    .A4(_1616_),
    .ZN(_2066_));
 NOR2_X1 _6263_ (.A1(_1324_),
    .A2(_1608_),
    .ZN(_2067_));
 AOI21_X1 _6264_ (.A(_2067_),
    .B1(_1607_),
    .B2(_1547_),
    .ZN(_2068_));
 NAND4_X1 _6265_ (.A1(\fir.p5[11] ),
    .A2(_1408_),
    .A3(_1544_),
    .A4(_1605_),
    .ZN(_2069_));
 AND3_X1 _6266_ (.A1(\fir.p5[11] ),
    .A2(_1513_),
    .A3(_1605_),
    .ZN(_2070_));
 NOR2_X1 _6267_ (.A1(_1551_),
    .A2(_1602_),
    .ZN(_2071_));
 INV_X1 _6268_ (.A(_1549_),
    .ZN(_2072_));
 AOI21_X1 _6269_ (.A(_2071_),
    .B1(_1603_),
    .B2(_2072_),
    .ZN(_2073_));
 NOR2_X1 _6270_ (.A1(_1556_),
    .A2(_1558_),
    .ZN(_2074_));
 INV_X1 _6271_ (.A(_1555_),
    .ZN(_2075_));
 AOI21_X1 _6272_ (.A(_2074_),
    .B1(_1559_),
    .B2(_2075_),
    .ZN(_2076_));
 OAI21_X1 _6273_ (.A(_1017_),
    .B1(_1040_),
    .B2(_0465_),
    .ZN(_2077_));
 OR2_X1 _6274_ (.A1(_1017_),
    .A2(_1040_),
    .ZN(_2078_));
 AND2_X1 _6275_ (.A1(_2077_),
    .A2(_2078_),
    .ZN(_2079_));
 NOR2_X1 _6276_ (.A1(_1566_),
    .A2(_1593_),
    .ZN(_2080_));
 NOR2_X1 _6277_ (.A1(_1563_),
    .A2(_1594_),
    .ZN(_2081_));
 NOR2_X1 _6278_ (.A1(_2080_),
    .A2(_2081_),
    .ZN(_2082_));
 NAND2_X1 _6279_ (.A1(\fir.p4[11] ),
    .A2(_1497_),
    .ZN(_2083_));
 MUX2_X1 _6280_ (.A(_0026_),
    .B(_2083_),
    .S(_1587_),
    .Z(_2084_));
 NAND2_X1 _6281_ (.A1(_1571_),
    .A2(_1585_),
    .ZN(_2085_));
 OAI21_X1 _6282_ (.A(_2085_),
    .B1(_1586_),
    .B2(_1569_),
    .ZN(_2086_));
 OAI21_X1 _6283_ (.A(_1582_),
    .B1(_1584_),
    .B2(_1368_),
    .ZN(_2087_));
 NAND2_X1 _6284_ (.A1(\fir.p2[11] ),
    .A2(_1578_),
    .ZN(_2088_));
 OAI21_X1 _6285_ (.A(_1248_),
    .B1(_1573_),
    .B2(_1577_),
    .ZN(_2089_));
 OAI211_X1 _6286_ (.A(_2088_),
    .B(_2089_),
    .C1(_1572_),
    .C2(_1578_),
    .ZN(_2090_));
 INV_X1 _6287_ (.A(_2090_),
    .ZN(_2091_));
 XNOR2_X1 _6288_ (.A(_2087_),
    .B(_2091_),
    .ZN(_2092_));
 XOR2_X1 _6289_ (.A(_2086_),
    .B(_2092_),
    .Z(_2093_));
 NOR2_X1 _6290_ (.A1(_0488_),
    .A2(_1587_),
    .ZN(_2094_));
 XNOR2_X1 _6291_ (.A(_2093_),
    .B(_2094_),
    .ZN(_2095_));
 XNOR2_X1 _6292_ (.A(_2084_),
    .B(_2095_),
    .ZN(_2096_));
 XNOR2_X1 _6293_ (.A(_1591_),
    .B(_2096_),
    .ZN(_2097_));
 MUX2_X1 _6294_ (.A(_1590_),
    .B(_0026_),
    .S(_1589_),
    .Z(_2098_));
 XOR2_X1 _6295_ (.A(_2097_),
    .B(_2098_),
    .Z(_2099_));
 XOR2_X1 _6296_ (.A(\fir.p4[11] ),
    .B(\fir.p3[11] ),
    .Z(_2100_));
 XOR2_X1 _6297_ (.A(_2099_),
    .B(_2100_),
    .Z(_2101_));
 XNOR2_X1 _6298_ (.A(_2082_),
    .B(_2101_),
    .ZN(_2102_));
 XNOR2_X1 _6299_ (.A(_2079_),
    .B(_2102_),
    .ZN(_2103_));
 NAND2_X1 _6300_ (.A1(_1560_),
    .A2(_1596_),
    .ZN(_2104_));
 OR2_X1 _6301_ (.A1(_1562_),
    .A2(_1595_),
    .ZN(_2105_));
 AOI21_X1 _6302_ (.A(_2103_),
    .B1(_2104_),
    .B2(_2105_),
    .ZN(_2106_));
 AND3_X1 _6303_ (.A1(_2105_),
    .A2(_2104_),
    .A3(_2103_),
    .ZN(_2107_));
 OR2_X1 _6304_ (.A1(_2106_),
    .A2(_2107_),
    .ZN(_2108_));
 XNOR2_X1 _6305_ (.A(_2076_),
    .B(_2108_),
    .ZN(_2109_));
 NAND2_X1 _6306_ (.A1(_1554_),
    .A2(_1601_),
    .ZN(_2110_));
 AOI21_X1 _6307_ (.A(_2109_),
    .B1(_2110_),
    .B2(_1599_),
    .ZN(_2111_));
 AND3_X1 _6308_ (.A1(_1599_),
    .A2(_2110_),
    .A3(_2109_),
    .ZN(_2112_));
 NOR2_X1 _6309_ (.A1(_2111_),
    .A2(_2112_),
    .ZN(_2113_));
 XNOR2_X1 _6310_ (.A(_2073_),
    .B(_2113_),
    .ZN(_2114_));
 OR2_X1 _6311_ (.A1(_0575_),
    .A2(_1604_),
    .ZN(_2115_));
 XNOR2_X1 _6312_ (.A(_2114_),
    .B(_2115_),
    .ZN(_2116_));
 XNOR2_X1 _6313_ (.A(_2070_),
    .B(_2116_),
    .ZN(_2117_));
 XOR2_X1 _6314_ (.A(_2069_),
    .B(_2117_),
    .Z(_2118_));
 XNOR2_X1 _6315_ (.A(\fir.p5[11] ),
    .B(_2118_),
    .ZN(_2119_));
 XNOR2_X1 _6316_ (.A(_2068_),
    .B(_2119_),
    .ZN(_2120_));
 NOR2_X1 _6317_ (.A1(_1542_),
    .A2(_1609_),
    .ZN(_2121_));
 AOI21_X1 _6318_ (.A(_1612_),
    .B1(_1542_),
    .B2(_1609_),
    .ZN(_2122_));
 AOI21_X1 _6319_ (.A(_2121_),
    .B1(_2122_),
    .B2(_1521_),
    .ZN(_2123_));
 XOR2_X1 _6320_ (.A(_2120_),
    .B(_2123_),
    .Z(_2124_));
 OAI21_X1 _6321_ (.A(\fir.p7[11] ),
    .B1(_1614_),
    .B2(_1615_),
    .ZN(_2125_));
 XOR2_X1 _6322_ (.A(_2124_),
    .B(_2125_),
    .Z(_2126_));
 XNOR2_X1 _6323_ (.A(_2066_),
    .B(_2126_),
    .ZN(_2127_));
 XNOR2_X1 _6324_ (.A(_1315_),
    .B(_2127_),
    .ZN(_2128_));
 XOR2_X1 _6325_ (.A(_2065_),
    .B(_2128_),
    .Z(_2129_));
 XNOR2_X1 _6326_ (.A(_1429_),
    .B(_2129_),
    .ZN(_2130_));
 XNOR2_X1 _6327_ (.A(_2062_),
    .B(_2130_),
    .ZN(_2131_));
 XOR2_X1 _6328_ (.A(_1537_),
    .B(_2131_),
    .Z(_2132_));
 XNOR2_X1 _6329_ (.A(_2059_),
    .B(_2132_),
    .ZN(_2133_));
 XOR2_X1 _6330_ (.A(_2057_),
    .B(_2133_),
    .Z(_2134_));
 AND2_X1 _6331_ (.A1(_1532_),
    .A2(_1627_),
    .ZN(_2135_));
 INV_X1 _6332_ (.A(_2135_),
    .ZN(_2136_));
 INV_X1 _6333_ (.A(_1628_),
    .ZN(_2137_));
 OAI21_X1 _6334_ (.A(_2136_),
    .B1(_2137_),
    .B2(_2038_),
    .ZN(_2138_));
 XNOR2_X1 _6335_ (.A(_2134_),
    .B(_2138_),
    .ZN(_2139_));
 OAI21_X1 _6336_ (.A(_2962_),
    .B1(_2056_),
    .B2(_2139_),
    .ZN(_2140_));
 AOI21_X1 _6337_ (.A(_2140_),
    .B1(_2139_),
    .B2(_2056_),
    .ZN(_0214_));
 AOI21_X1 _6338_ (.A(_2039_),
    .B1(_2053_),
    .B2(_2055_),
    .ZN(_2141_));
 NAND2_X1 _6339_ (.A1(_2962_),
    .A2(_2056_),
    .ZN(_2142_));
 NOR2_X1 _6340_ (.A1(_2141_),
    .A2(_2142_),
    .ZN(_0213_));
 OAI21_X1 _6341_ (.A(_2962_),
    .B1(_2053_),
    .B2(_2055_),
    .ZN(_2143_));
 AOI21_X1 _6342_ (.A(_2143_),
    .B1(_2055_),
    .B2(_2053_),
    .ZN(_0212_));
 NOR2_X1 _6343_ (.A1(_2040_),
    .A2(_2052_),
    .ZN(_2144_));
 NOR3_X1 _6344_ (.A1(rst),
    .A2(_2053_),
    .A3(_2144_),
    .ZN(_0211_));
 NOR2_X1 _6345_ (.A1(_2041_),
    .A2(_2051_),
    .ZN(_2145_));
 NOR3_X1 _6346_ (.A1(rst),
    .A2(_2052_),
    .A3(_2145_),
    .ZN(_0210_));
 NOR2_X1 _6347_ (.A1(_2042_),
    .A2(_2050_),
    .ZN(_2146_));
 NOR3_X1 _6348_ (.A1(rst),
    .A2(_2051_),
    .A3(_2146_),
    .ZN(_0209_));
 AND2_X1 _6349_ (.A1(_2048_),
    .A2(_2049_),
    .ZN(_2147_));
 NOR3_X1 _6350_ (.A1(rst),
    .A2(_2050_),
    .A3(_2147_),
    .ZN(_0208_));
 OAI21_X1 _6351_ (.A(_2962_),
    .B1(_2043_),
    .B2(_2047_),
    .ZN(_2148_));
 AOI21_X1 _6352_ (.A(_2148_),
    .B1(_2047_),
    .B2(_2043_),
    .ZN(_0207_));
 AOI21_X1 _6353_ (.A(_2046_),
    .B1(_2045_),
    .B2(_2044_),
    .ZN(_2149_));
 NOR3_X1 _6354_ (.A1(rst),
    .A2(_2047_),
    .A3(_2149_),
    .ZN(_0206_));
 INV_X1 _6355_ (.A(_2132_),
    .ZN(_2150_));
 NOR2_X1 _6356_ (.A1(_2059_),
    .A2(_2150_),
    .ZN(_2151_));
 INV_X1 _6357_ (.A(_2130_),
    .ZN(_2152_));
 NOR2_X1 _6358_ (.A1(_2062_),
    .A2(_2152_),
    .ZN(_2153_));
 AOI21_X1 _6359_ (.A(_2153_),
    .B1(_2131_),
    .B2(_1537_),
    .ZN(_2154_));
 NAND2_X1 _6360_ (.A1(_2061_),
    .A2(_2129_),
    .ZN(_2155_));
 OAI21_X1 _6361_ (.A(_2155_),
    .B1(_2128_),
    .B2(_2065_),
    .ZN(_2156_));
 AND2_X1 _6362_ (.A1(_2066_),
    .A2(_2126_),
    .ZN(_2157_));
 NOR2_X1 _6363_ (.A1(_1315_),
    .A2(_2127_),
    .ZN(_2158_));
 NOR2_X1 _6364_ (.A1(_2157_),
    .A2(_2158_),
    .ZN(_2159_));
 NAND3_X1 _6365_ (.A1(\fir.p7[11] ),
    .A2(_1616_),
    .A3(_2124_),
    .ZN(_2160_));
 NOR2_X1 _6366_ (.A1(_2068_),
    .A2(_2119_),
    .ZN(_2161_));
 AOI211_X1 _6367_ (.A(_2121_),
    .B(_2120_),
    .C1(_2122_),
    .C2(_1521_),
    .ZN(_2162_));
 NAND2_X1 _6368_ (.A1(_2069_),
    .A2(_2117_),
    .ZN(_2163_));
 NAND2_X1 _6369_ (.A1(\fir.p5[11] ),
    .A2(_2163_),
    .ZN(_2164_));
 AND2_X1 _6370_ (.A1(_2070_),
    .A2(_2116_),
    .ZN(_2165_));
 NOR2_X1 _6371_ (.A1(_2114_),
    .A2(_2115_),
    .ZN(_2166_));
 NOR2_X1 _6372_ (.A1(_2076_),
    .A2(_2108_),
    .ZN(_2167_));
 NOR2_X1 _6373_ (.A1(_2106_),
    .A2(_2167_),
    .ZN(_2168_));
 INV_X1 _6374_ (.A(_2078_),
    .ZN(_2169_));
 NOR2_X1 _6375_ (.A1(\fir.p4[11] ),
    .A2(_0465_),
    .ZN(_2170_));
 MUX2_X1 _6376_ (.A(_0026_),
    .B(_2084_),
    .S(_2095_),
    .Z(_2171_));
 NAND2_X1 _6377_ (.A1(_2087_),
    .A2(_2091_),
    .ZN(_2172_));
 INV_X1 _6378_ (.A(_2086_),
    .ZN(_2173_));
 OAI211_X1 _6379_ (.A(_2089_),
    .B(_2172_),
    .C1(_2092_),
    .C2(_2173_),
    .ZN(_2174_));
 NAND2_X1 _6380_ (.A1(\fir.p4[11] ),
    .A2(_2093_),
    .ZN(_2175_));
 XOR2_X1 _6381_ (.A(_2174_),
    .B(_2175_),
    .Z(_2176_));
 NAND2_X1 _6382_ (.A1(\fir.p4[11] ),
    .A2(_1587_),
    .ZN(_2177_));
 INV_X1 _6383_ (.A(_2093_),
    .ZN(_2178_));
 NAND2_X1 _6384_ (.A1(_2177_),
    .A2(_2178_),
    .ZN(_2179_));
 OAI21_X1 _6385_ (.A(_0026_),
    .B1(_2177_),
    .B2(_2093_),
    .ZN(_2180_));
 NAND2_X1 _6386_ (.A1(_2179_),
    .A2(_2180_),
    .ZN(_2181_));
 XNOR2_X1 _6387_ (.A(_1591_),
    .B(_2181_),
    .ZN(_2182_));
 XNOR2_X1 _6388_ (.A(_2176_),
    .B(_2182_),
    .ZN(_2183_));
 XOR2_X1 _6389_ (.A(_2171_),
    .B(_2183_),
    .Z(_2184_));
 XOR2_X1 _6390_ (.A(_2100_),
    .B(_2184_),
    .Z(_2185_));
 AND2_X1 _6391_ (.A1(_2099_),
    .A2(_2100_),
    .ZN(_2186_));
 NOR2_X1 _6392_ (.A1(_2097_),
    .A2(_2098_),
    .ZN(_2187_));
 OAI21_X1 _6393_ (.A(_2185_),
    .B1(_2186_),
    .B2(_2187_),
    .ZN(_2188_));
 OR3_X1 _6394_ (.A1(_2187_),
    .A2(_2186_),
    .A3(_2185_),
    .ZN(_2189_));
 AND2_X1 _6395_ (.A1(_2188_),
    .A2(_2189_),
    .ZN(_2190_));
 XNOR2_X1 _6396_ (.A(_2170_),
    .B(_2190_),
    .ZN(_2191_));
 NAND2_X1 _6397_ (.A1(_2079_),
    .A2(_2102_),
    .ZN(_2192_));
 OAI21_X1 _6398_ (.A(_2101_),
    .B1(_2081_),
    .B2(_2080_),
    .ZN(_2193_));
 AOI21_X1 _6399_ (.A(_2191_),
    .B1(_2192_),
    .B2(_2193_),
    .ZN(_2194_));
 AND3_X1 _6400_ (.A1(_2193_),
    .A2(_2192_),
    .A3(_2191_),
    .ZN(_2195_));
 NOR2_X1 _6401_ (.A1(_2194_),
    .A2(_2195_),
    .ZN(_2196_));
 XNOR2_X1 _6402_ (.A(_2169_),
    .B(_2196_),
    .ZN(_2197_));
 XOR2_X1 _6403_ (.A(_2168_),
    .B(_2197_),
    .Z(_2198_));
 INV_X1 _6404_ (.A(_2113_),
    .ZN(_2199_));
 NOR2_X1 _6405_ (.A1(_2073_),
    .A2(_2199_),
    .ZN(_2200_));
 OAI21_X1 _6406_ (.A(_2198_),
    .B1(_2200_),
    .B2(_2111_),
    .ZN(_2201_));
 OR3_X1 _6407_ (.A1(_2111_),
    .A2(_2200_),
    .A3(_2198_),
    .ZN(_2202_));
 AND2_X1 _6408_ (.A1(_2201_),
    .A2(_2202_),
    .ZN(_2203_));
 XOR2_X1 _6409_ (.A(_2166_),
    .B(_2203_),
    .Z(_2204_));
 OR2_X1 _6410_ (.A1(_2165_),
    .A2(_2204_),
    .ZN(_2205_));
 NAND2_X1 _6411_ (.A1(_2165_),
    .A2(_2204_),
    .ZN(_2206_));
 NAND3_X1 _6412_ (.A1(\fir.p5[11] ),
    .A2(_2205_),
    .A3(_2206_),
    .ZN(_2207_));
 OAI21_X1 _6413_ (.A(_2207_),
    .B1(_2203_),
    .B2(\fir.p5[11] ),
    .ZN(_2208_));
 XOR2_X1 _6414_ (.A(_2164_),
    .B(_2208_),
    .Z(_2209_));
 OR3_X1 _6415_ (.A1(_2161_),
    .A2(_2162_),
    .A3(_2209_),
    .ZN(_2210_));
 OAI21_X1 _6416_ (.A(_2209_),
    .B1(_2162_),
    .B2(_2161_),
    .ZN(_2211_));
 AND2_X1 _6417_ (.A1(_2210_),
    .A2(_2211_),
    .ZN(_2212_));
 XOR2_X1 _6418_ (.A(_2160_),
    .B(_2212_),
    .Z(_2213_));
 XOR2_X1 _6419_ (.A(_1315_),
    .B(_2213_),
    .Z(_2214_));
 XNOR2_X1 _6420_ (.A(_2159_),
    .B(_2214_),
    .ZN(_2215_));
 XNOR2_X1 _6421_ (.A(_1429_),
    .B(_2215_),
    .ZN(_2216_));
 XOR2_X1 _6422_ (.A(_2156_),
    .B(_2216_),
    .Z(_2217_));
 XNOR2_X1 _6423_ (.A(_1537_),
    .B(_2217_),
    .ZN(_2218_));
 XOR2_X1 _6424_ (.A(_2154_),
    .B(_2218_),
    .Z(_2219_));
 AND2_X1 _6425_ (.A1(_2151_),
    .A2(_2219_),
    .ZN(_2220_));
 XOR2_X1 _6426_ (.A(_2151_),
    .B(_2219_),
    .Z(_2221_));
 AND2_X1 _6427_ (.A1(_2057_),
    .A2(_2133_),
    .ZN(_2222_));
 AOI21_X1 _6428_ (.A(_2222_),
    .B1(_2134_),
    .B2(_2135_),
    .ZN(_2223_));
 NAND4_X1 _6429_ (.A1(_1628_),
    .A2(_2037_),
    .A3(_1697_),
    .A4(_2134_),
    .ZN(_2224_));
 NAND2_X1 _6430_ (.A1(_1628_),
    .A2(_2134_),
    .ZN(_2225_));
 AOI21_X1 _6431_ (.A(_1657_),
    .B1(_1694_),
    .B2(_1695_),
    .ZN(_2226_));
 OAI211_X1 _6432_ (.A(_2223_),
    .B(_2224_),
    .C1(_2225_),
    .C2(_2226_),
    .ZN(_2227_));
 AOI21_X1 _6433_ (.A(_2220_),
    .B1(_2221_),
    .B2(_2227_),
    .ZN(_2228_));
 NOR2_X1 _6434_ (.A1(_2154_),
    .A2(_2218_),
    .ZN(_2229_));
 AND2_X1 _6435_ (.A1(_2156_),
    .A2(_2216_),
    .ZN(_2230_));
 AOI21_X1 _6436_ (.A(_2230_),
    .B1(_2217_),
    .B2(_1537_),
    .ZN(_2231_));
 OAI21_X1 _6437_ (.A(_2214_),
    .B1(_2158_),
    .B2(_2157_),
    .ZN(_2232_));
 INV_X1 _6438_ (.A(_2215_),
    .ZN(_2233_));
 OAI21_X1 _6439_ (.A(_2232_),
    .B1(_2233_),
    .B2(_1429_),
    .ZN(_2234_));
 NAND2_X1 _6440_ (.A1(\fir.p7[11] ),
    .A2(_2124_),
    .ZN(_2235_));
 OR3_X1 _6441_ (.A1(_1616_),
    .A2(_2212_),
    .A3(_2235_),
    .ZN(_2236_));
 OAI21_X1 _6442_ (.A(_2236_),
    .B1(_2213_),
    .B2(_1315_),
    .ZN(_2237_));
 OAI21_X1 _6443_ (.A(_2211_),
    .B1(_2208_),
    .B2(_2164_),
    .ZN(_2238_));
 NAND2_X1 _6444_ (.A1(_2206_),
    .A2(_2207_),
    .ZN(_2239_));
 OAI21_X1 _6445_ (.A(_2201_),
    .B1(_2197_),
    .B2(_2168_),
    .ZN(_2240_));
 AOI21_X1 _6446_ (.A(_2194_),
    .B1(_2196_),
    .B2(_2169_),
    .ZN(_2241_));
 INV_X1 _6447_ (.A(_2188_),
    .ZN(_2242_));
 AOI21_X1 _6448_ (.A(_2242_),
    .B1(_2190_),
    .B2(_2170_),
    .ZN(_2243_));
 NOR2_X1 _6449_ (.A1(_2171_),
    .A2(_2183_),
    .ZN(_2244_));
 AOI21_X1 _6450_ (.A(_2244_),
    .B1(_2184_),
    .B2(_2100_),
    .ZN(_2245_));
 OAI211_X1 _6451_ (.A(_2176_),
    .B(_2180_),
    .C1(_2181_),
    .C2(_0026_),
    .ZN(_2246_));
 AOI21_X1 _6452_ (.A(_2174_),
    .B1(_2178_),
    .B2(\fir.p4[11] ),
    .ZN(_2247_));
 XNOR2_X1 _6453_ (.A(_2246_),
    .B(_2247_),
    .ZN(_2248_));
 XOR2_X1 _6454_ (.A(_2245_),
    .B(_2248_),
    .Z(_2249_));
 XNOR2_X1 _6455_ (.A(_2243_),
    .B(_2249_),
    .ZN(_2250_));
 XNOR2_X1 _6456_ (.A(_2241_),
    .B(_2250_),
    .ZN(_2251_));
 XNOR2_X1 _6457_ (.A(_2240_),
    .B(_2251_),
    .ZN(_2252_));
 NOR3_X1 _6458_ (.A1(_1604_),
    .A2(_2114_),
    .A3(_2203_),
    .ZN(_2253_));
 NOR2_X1 _6459_ (.A1(_0575_),
    .A2(_2253_),
    .ZN(_2254_));
 XNOR2_X1 _6460_ (.A(_2252_),
    .B(_2254_),
    .ZN(_2255_));
 XNOR2_X1 _6461_ (.A(_2239_),
    .B(_2255_),
    .ZN(_2256_));
 XNOR2_X1 _6462_ (.A(_2238_),
    .B(_2256_),
    .ZN(_2257_));
 OAI21_X1 _6463_ (.A(\fir.p7[11] ),
    .B1(_2212_),
    .B2(_2235_),
    .ZN(_2258_));
 XNOR2_X1 _6464_ (.A(_2257_),
    .B(_2258_),
    .ZN(_2259_));
 XNOR2_X1 _6465_ (.A(_2237_),
    .B(_2259_),
    .ZN(_2260_));
 XNOR2_X1 _6466_ (.A(_2234_),
    .B(_2260_),
    .ZN(_2261_));
 XNOR2_X1 _6467_ (.A(_2231_),
    .B(_2261_),
    .ZN(_2262_));
 XNOR2_X1 _6468_ (.A(_2229_),
    .B(_2262_),
    .ZN(_2263_));
 XNOR2_X1 _6469_ (.A(_2228_),
    .B(_2263_),
    .ZN(_2264_));
 XNOR2_X1 _6470_ (.A(_2221_),
    .B(_2227_),
    .ZN(_2265_));
 NOR3_X1 _6471_ (.A1(_2056_),
    .A2(_2139_),
    .A3(_2265_),
    .ZN(_2266_));
 OAI21_X1 _6472_ (.A(_2962_),
    .B1(_2264_),
    .B2(_2266_),
    .ZN(_2267_));
 AOI21_X1 _6473_ (.A(_2267_),
    .B1(_2266_),
    .B2(_2264_),
    .ZN(_0205_));
 OAI21_X1 _6474_ (.A(_2265_),
    .B1(_2139_),
    .B2(_2056_),
    .ZN(_2268_));
 NAND2_X1 _6475_ (.A1(_2962_),
    .A2(_2268_),
    .ZN(_2269_));
 NOR2_X1 _6476_ (.A1(_2266_),
    .A2(_2269_),
    .ZN(_0204_));
 OAI21_X1 _6477_ (.A(_2962_),
    .B1(_2044_),
    .B2(_2045_),
    .ZN(_2270_));
 AOI21_X1 _6478_ (.A(_2270_),
    .B1(_2045_),
    .B2(_2044_),
    .ZN(_0203_));
 AND2_X1 _6479_ (.A1(_2962_),
    .A2(net149),
    .ZN(_0202_));
 AND2_X1 _6480_ (.A1(_2962_),
    .A2(net147),
    .ZN(_0201_));
 AND2_X1 _6481_ (.A1(_2962_),
    .A2(net143),
    .ZN(_0200_));
 AND2_X1 _6482_ (.A1(_2962_),
    .A2(net223),
    .ZN(_0199_));
 AND2_X1 _6483_ (.A1(_2962_),
    .A2(net263),
    .ZN(_0198_));
 AND2_X1 _6484_ (.A1(_2962_),
    .A2(net249),
    .ZN(_0197_));
 AND2_X1 _6485_ (.A1(_2962_),
    .A2(net259),
    .ZN(_0196_));
 AND2_X1 _6486_ (.A1(_2962_),
    .A2(net215),
    .ZN(_0195_));
 NOR2_X1 _6487_ (.A1(rst),
    .A2(net214),
    .ZN(_0194_));
 NOR2_X1 _6488_ (.A1(rst),
    .A2(net170),
    .ZN(_0193_));
 AND2_X1 _6489_ (.A1(_2962_),
    .A2(net137),
    .ZN(_0192_));
 NOR2_X1 _6490_ (.A1(rst),
    .A2(net121),
    .ZN(_0191_));
 AND2_X1 _6491_ (.A1(_2962_),
    .A2(net199),
    .ZN(_0190_));
 AND2_X1 _6492_ (.A1(_2962_),
    .A2(net181),
    .ZN(_0189_));
 AND2_X1 _6493_ (.A1(_2962_),
    .A2(net197),
    .ZN(_0188_));
 NOR2_X1 _6494_ (.A1(rst),
    .A2(net186),
    .ZN(_0187_));
 AND2_X1 _6495_ (.A1(_2962_),
    .A2(net175),
    .ZN(_0186_));
 AND2_X1 _6496_ (.A1(_2962_),
    .A2(net179),
    .ZN(_0185_));
 AND2_X1 _6497_ (.A1(_2962_),
    .A2(net171),
    .ZN(_0184_));
 AND2_X1 _6498_ (.A1(_2962_),
    .A2(net189),
    .ZN(_0183_));
 AND2_X1 _6499_ (.A1(_2962_),
    .A2(net159),
    .ZN(_0182_));
 NOR2_X1 _6500_ (.A1(rst),
    .A2(_0575_),
    .ZN(_0181_));
 NOR2_X1 _6501_ (.A1(rst),
    .A2(net230),
    .ZN(_0180_));
 AND2_X1 _6502_ (.A1(_2962_),
    .A2(net183),
    .ZN(_0179_));
 AND2_X1 _6503_ (.A1(_2962_),
    .A2(net261),
    .ZN(_0178_));
 NOR2_X1 _6504_ (.A1(rst),
    .A2(net268),
    .ZN(_0177_));
 AND2_X1 _6505_ (.A1(_2962_),
    .A2(net253),
    .ZN(_0176_));
 AND2_X1 _6506_ (.A1(_2962_),
    .A2(net257),
    .ZN(_0175_));
 AND2_X1 _6507_ (.A1(_2962_),
    .A2(net255),
    .ZN(_0174_));
 AND2_X1 _6508_ (.A1(_2962_),
    .A2(net251),
    .ZN(_0173_));
 AND2_X1 _6509_ (.A1(_2962_),
    .A2(net237),
    .ZN(_0172_));
 AND2_X1 _6510_ (.A1(_2962_),
    .A2(net239),
    .ZN(_0171_));
 NOR2_X1 _6511_ (.A1(rst),
    .A2(net280),
    .ZN(_0170_));
 NOR2_X1 _6512_ (.A1(rst),
    .A2(_0488_),
    .ZN(_0169_));
 AND2_X1 _6513_ (.A1(_2962_),
    .A2(net241),
    .ZN(_0168_));
 AND2_X1 _6514_ (.A1(_2962_),
    .A2(net275),
    .ZN(_0167_));
 AND2_X1 _6515_ (.A1(_2962_),
    .A2(net271),
    .ZN(_0166_));
 AND2_X1 _6516_ (.A1(_2962_),
    .A2(net219),
    .ZN(_0165_));
 AND2_X1 _6517_ (.A1(_2962_),
    .A2(net221),
    .ZN(_0164_));
 AND2_X1 _6518_ (.A1(_2962_),
    .A2(net217),
    .ZN(_0163_));
 AND2_X1 _6519_ (.A1(_2962_),
    .A2(net245),
    .ZN(_0162_));
 AND2_X1 _6520_ (.A1(_2962_),
    .A2(net211),
    .ZN(_0161_));
 AND2_X1 _6521_ (.A1(_2962_),
    .A2(net247),
    .ZN(_0160_));
 AND2_X1 _6522_ (.A1(_2962_),
    .A2(net209),
    .ZN(_0159_));
 AND2_X1 _6523_ (.A1(_2962_),
    .A2(net269),
    .ZN(_0158_));
 NOR2_X1 _6524_ (.A1(rst),
    .A2(_0465_),
    .ZN(_0157_));
 AND2_X1 _6525_ (.A1(_2962_),
    .A2(net273),
    .ZN(_0156_));
 AND2_X1 _6526_ (.A1(_2962_),
    .A2(net277),
    .ZN(_0155_));
 AND2_X1 _6527_ (.A1(_2962_),
    .A2(net193),
    .ZN(_0154_));
 AND2_X1 _6528_ (.A1(_2962_),
    .A2(net165),
    .ZN(_0153_));
 AND2_X1 _6529_ (.A1(_2962_),
    .A2(net135),
    .ZN(_0152_));
 AND2_X1 _6530_ (.A1(_2962_),
    .A2(net133),
    .ZN(_0151_));
 AND2_X1 _6531_ (.A1(_2962_),
    .A2(net163),
    .ZN(_0150_));
 AND2_X1 _6532_ (.A1(_2962_),
    .A2(net191),
    .ZN(_0149_));
 AND2_X1 _6533_ (.A1(_2962_),
    .A2(net145),
    .ZN(_0148_));
 AND2_X1 _6534_ (.A1(_2962_),
    .A2(net139),
    .ZN(_0147_));
 AND2_X1 _6535_ (.A1(_2962_),
    .A2(net167),
    .ZN(_0146_));
 NOR2_X1 _6536_ (.A1(rst),
    .A2(_1248_),
    .ZN(_0145_));
 AND2_X1 _6537_ (.A1(_2962_),
    .A2(net195),
    .ZN(_0144_));
 AND2_X1 _6538_ (.A1(_2962_),
    .A2(net187),
    .ZN(_0143_));
 AND2_X1 _6539_ (.A1(_2962_),
    .A2(net201),
    .ZN(_0142_));
 AND2_X1 _6540_ (.A1(_2962_),
    .A2(net243),
    .ZN(_0141_));
 AND2_X1 _6541_ (.A1(_2962_),
    .A2(net231),
    .ZN(_0140_));
 AND2_X1 _6542_ (.A1(_2962_),
    .A2(net151),
    .ZN(_0139_));
 AND2_X1 _6543_ (.A1(_2962_),
    .A2(net157),
    .ZN(_0138_));
 AND2_X1 _6544_ (.A1(_2962_),
    .A2(net131),
    .ZN(_0137_));
 AND2_X1 _6545_ (.A1(_2962_),
    .A2(net141),
    .ZN(_0136_));
 AND2_X1 _6546_ (.A1(_2962_),
    .A2(net173),
    .ZN(_0135_));
 AND2_X1 _6547_ (.A1(_2962_),
    .A2(net118),
    .ZN(_0134_));
 NOR2_X1 _6548_ (.A1(rst),
    .A2(net266),
    .ZN(_0133_));
 AND2_X1 _6549_ (.A1(_2962_),
    .A2(net205),
    .ZN(_0132_));
 AND2_X1 _6550_ (.A1(_2962_),
    .A2(net113),
    .ZN(_0131_));
 AND2_X1 _6551_ (.A1(_2962_),
    .A2(net126),
    .ZN(_0130_));
 AND2_X1 _6552_ (.A1(_2962_),
    .A2(net227),
    .ZN(_0129_));
 AND2_X1 _6553_ (.A1(_2962_),
    .A2(net225),
    .ZN(_0128_));
 AND2_X1 _6554_ (.A1(_2962_),
    .A2(net235),
    .ZN(_0127_));
 AND2_X1 _6555_ (.A1(_2962_),
    .A2(net207),
    .ZN(_0126_));
 AND2_X1 _6556_ (.A1(_2962_),
    .A2(net233),
    .ZN(_0125_));
 AND2_X1 _6557_ (.A1(_2962_),
    .A2(net203),
    .ZN(_0124_));
 AND2_X1 _6558_ (.A1(_2962_),
    .A2(net177),
    .ZN(_0123_));
 AND2_X1 _6559_ (.A1(_2962_),
    .A2(net161),
    .ZN(_0122_));
 NOR2_X1 _6560_ (.A1(rst),
    .A2(net129),
    .ZN(_0121_));
 AND2_X1 _6561_ (.A1(_2962_),
    .A2(net155),
    .ZN(_0120_));
 AND2_X1 _6562_ (.A1(_2962_),
    .A2(net153),
    .ZN(_0119_));
 AND2_X1 _6563_ (.A1(_2962_),
    .A2(net390),
    .ZN(_0118_));
 AND2_X1 _6564_ (.A1(_2962_),
    .A2(net320),
    .ZN(_0117_));
 AND2_X1 _6565_ (.A1(_2962_),
    .A2(net358),
    .ZN(_0116_));
 AND2_X1 _6566_ (.A1(_2962_),
    .A2(net340),
    .ZN(_0115_));
 AND2_X1 _6567_ (.A1(_2962_),
    .A2(net396),
    .ZN(_0114_));
 AND2_X1 _6568_ (.A1(_2962_),
    .A2(net394),
    .ZN(_0113_));
 AND2_X1 _6569_ (.A1(_2962_),
    .A2(net370),
    .ZN(_0112_));
 AND2_X1 _6570_ (.A1(_2962_),
    .A2(net344),
    .ZN(_0111_));
 AND2_X1 _6571_ (.A1(_2962_),
    .A2(net342),
    .ZN(_0110_));
 AND2_X1 _6572_ (.A1(_2962_),
    .A2(net386),
    .ZN(_0109_));
 AND2_X1 _6573_ (.A1(_2962_),
    .A2(net382),
    .ZN(_0108_));
 AND2_X1 _6574_ (.A1(_2962_),
    .A2(net109),
    .ZN(_0107_));
 AND2_X1 _6575_ (.A1(_2962_),
    .A2(net310),
    .ZN(_0106_));
 AND2_X1 _6576_ (.A1(_2962_),
    .A2(net338),
    .ZN(_0105_));
 AND2_X1 _6577_ (.A1(_2962_),
    .A2(net378),
    .ZN(_0104_));
 AND2_X1 _6578_ (.A1(_2962_),
    .A2(net368),
    .ZN(_0103_));
 AND2_X1 _6579_ (.A1(_2962_),
    .A2(net366),
    .ZN(_0102_));
 AND2_X1 _6580_ (.A1(_2962_),
    .A2(net374),
    .ZN(_0101_));
 AND2_X1 _6581_ (.A1(_2962_),
    .A2(net372),
    .ZN(_0100_));
 AND2_X1 _6582_ (.A1(_2962_),
    .A2(net380),
    .ZN(_0099_));
 AND2_X1 _6583_ (.A1(_2962_),
    .A2(net362),
    .ZN(_0098_));
 AND2_X1 _6584_ (.A1(_2962_),
    .A2(net376),
    .ZN(_0097_));
 AND2_X1 _6585_ (.A1(_2962_),
    .A2(net364),
    .ZN(_0096_));
 AND2_X1 _6586_ (.A1(_2962_),
    .A2(net322),
    .ZN(_0095_));
 AND2_X1 _6587_ (.A1(_2962_),
    .A2(net334),
    .ZN(_0094_));
 AND2_X1 _6588_ (.A1(_2962_),
    .A2(net332),
    .ZN(_0093_));
 AND2_X1 _6589_ (.A1(_2962_),
    .A2(net302),
    .ZN(_0092_));
 AND2_X1 _6590_ (.A1(_2962_),
    .A2(net304),
    .ZN(_0091_));
 AND2_X1 _6591_ (.A1(_2962_),
    .A2(net346),
    .ZN(_0090_));
 AND2_X1 _6592_ (.A1(_2962_),
    .A2(net354),
    .ZN(_0089_));
 AND2_X1 _6593_ (.A1(_2962_),
    .A2(net360),
    .ZN(_0088_));
 AND2_X1 _6594_ (.A1(_2962_),
    .A2(net324),
    .ZN(_0087_));
 AND2_X1 _6595_ (.A1(_2962_),
    .A2(net356),
    .ZN(_0086_));
 AND2_X1 _6596_ (.A1(_2962_),
    .A2(net348),
    .ZN(_0085_));
 AND2_X1 _6597_ (.A1(_2962_),
    .A2(net326),
    .ZN(_0084_));
 AND2_X1 _6598_ (.A1(_2962_),
    .A2(net336),
    .ZN(_0083_));
 AND2_X1 _6599_ (.A1(_2962_),
    .A2(net314),
    .ZN(_0082_));
 AND2_X1 _6600_ (.A1(_2962_),
    .A2(net306),
    .ZN(_0081_));
 AND2_X1 _6601_ (.A1(_2962_),
    .A2(net308),
    .ZN(_0080_));
 AND2_X1 _6602_ (.A1(_2962_),
    .A2(net312),
    .ZN(_0079_));
 AND2_X1 _6603_ (.A1(_2962_),
    .A2(net330),
    .ZN(_0078_));
 AND2_X1 _6604_ (.A1(_2962_),
    .A2(net316),
    .ZN(_0077_));
 AND2_X1 _6605_ (.A1(_2962_),
    .A2(net318),
    .ZN(_0076_));
 AND2_X1 _6606_ (.A1(_2962_),
    .A2(net328),
    .ZN(_0075_));
 AND2_X1 _6607_ (.A1(_2962_),
    .A2(net350),
    .ZN(_0074_));
 INV_X1 _6608_ (.A(net290),
    .ZN(_2271_));
 NOR2_X1 _6609_ (.A1(rst),
    .A2(_2271_),
    .ZN(_0073_));
 INV_X1 _6610_ (.A(net288),
    .ZN(_2272_));
 NOR2_X1 _6611_ (.A1(rst),
    .A2(_2272_),
    .ZN(_0072_));
 INV_X1 _6612_ (.A(net284),
    .ZN(_2273_));
 NOR2_X1 _6613_ (.A1(rst),
    .A2(_2273_),
    .ZN(_0071_));
 INV_X1 _6614_ (.A(net281),
    .ZN(_2274_));
 NOR2_X1 _6615_ (.A1(rst),
    .A2(net282),
    .ZN(_0070_));
 AND2_X1 _6616_ (.A1(_2962_),
    .A2(net289),
    .ZN(_0069_));
 INV_X1 _6617_ (.A(net283),
    .ZN(_2275_));
 NOR2_X1 _6618_ (.A1(rst),
    .A2(_2275_),
    .ZN(_0068_));
 INV_X1 _6619_ (.A(net123),
    .ZN(_2276_));
 NOR2_X1 _6620_ (.A1(rst),
    .A2(net124),
    .ZN(_0067_));
 INV_X1 _6621_ (.A(net449),
    .ZN(_2277_));
 NOR2_X1 _6622_ (.A1(rst),
    .A2(_2277_),
    .ZN(_0066_));
 INV_X1 _6623_ (.A(net285),
    .ZN(_2278_));
 NOR2_X1 _6624_ (.A1(rst),
    .A2(_2278_),
    .ZN(_0065_));
 INV_X1 _6625_ (.A(net115),
    .ZN(_2279_));
 NOR2_X1 _6626_ (.A1(rst),
    .A2(net116),
    .ZN(_0064_));
 INV_X1 _6627_ (.A(net287),
    .ZN(_2280_));
 NOR2_X1 _6628_ (.A1(rst),
    .A2(_2280_),
    .ZN(_0063_));
 AND2_X1 _6629_ (.A1(_2962_),
    .A2(net292),
    .ZN(_0062_));
 AND2_X1 _6630_ (.A1(_2962_),
    .A2(net398),
    .ZN(_0061_));
 AND2_X1 _6631_ (.A1(_2962_),
    .A2(net392),
    .ZN(_0060_));
 AND2_X1 _6632_ (.A1(_2962_),
    .A2(net298),
    .ZN(_0059_));
 AND2_X1 _6633_ (.A1(_2962_),
    .A2(net300),
    .ZN(_0058_));
 AND2_X1 _6634_ (.A1(_2962_),
    .A2(net400),
    .ZN(_0057_));
 AND2_X1 _6635_ (.A1(_2962_),
    .A2(net352),
    .ZN(_0056_));
 AND2_X1 _6636_ (.A1(_2962_),
    .A2(net294),
    .ZN(_0055_));
 AND2_X1 _6637_ (.A1(_2962_),
    .A2(net388),
    .ZN(_0054_));
 AND2_X1 _6638_ (.A1(_2962_),
    .A2(net296),
    .ZN(_0053_));
 AND2_X1 _6639_ (.A1(_2962_),
    .A2(net384),
    .ZN(_0052_));
 NOR2_X1 _6640_ (.A1(_2273_),
    .A2(\aso.z4[7] ),
    .ZN(_2281_));
 XOR2_X1 _6641_ (.A(\aso.z0[6] ),
    .B(\aso.z4[6] ),
    .Z(_2282_));
 XOR2_X1 _6642_ (.A(\aso.z0[5] ),
    .B(\aso.z4[5] ),
    .Z(_2283_));
 NOR2_X1 _6643_ (.A1(_2275_),
    .A2(\aso.z4[4] ),
    .ZN(_2284_));
 OR2_X1 _6644_ (.A1(_2276_),
    .A2(\aso.z4[3] ),
    .ZN(_2285_));
 XOR2_X1 _6645_ (.A(\aso.z0[3] ),
    .B(\aso.z4[3] ),
    .Z(_2286_));
 NOR2_X1 _6646_ (.A1(_2277_),
    .A2(\aso.z4[2] ),
    .ZN(_2287_));
 NAND2_X1 _6647_ (.A1(_2280_),
    .A2(\aso.z4[0] ),
    .ZN(_2288_));
 XNOR2_X1 _6648_ (.A(\aso.z0[1] ),
    .B(\aso.z4[1] ),
    .ZN(_2289_));
 NAND2_X1 _6649_ (.A1(_2288_),
    .A2(_2289_),
    .ZN(_2290_));
 OAI21_X1 _6650_ (.A(_2290_),
    .B1(\aso.z4[1] ),
    .B2(_2278_),
    .ZN(_2291_));
 XNOR2_X1 _6651_ (.A(\aso.z0[2] ),
    .B(\aso.z4[2] ),
    .ZN(_2292_));
 AOI21_X1 _6652_ (.A(_2287_),
    .B1(_2291_),
    .B2(_2292_),
    .ZN(_2293_));
 OAI21_X1 _6653_ (.A(_2285_),
    .B1(_2286_),
    .B2(_2293_),
    .ZN(_2294_));
 XNOR2_X1 _6654_ (.A(\aso.z0[4] ),
    .B(\aso.z4[4] ),
    .ZN(_2295_));
 AOI21_X1 _6655_ (.A(_2284_),
    .B1(_2294_),
    .B2(_2295_),
    .ZN(_2296_));
 NOR2_X1 _6656_ (.A1(_2283_),
    .A2(_2296_),
    .ZN(_2297_));
 INV_X1 _6657_ (.A(\aso.z4[5] ),
    .ZN(_2298_));
 AOI21_X1 _6658_ (.A(_2297_),
    .B1(_2298_),
    .B2(\aso.z0[5] ),
    .ZN(_2299_));
 NOR2_X1 _6659_ (.A1(_2282_),
    .A2(_2299_),
    .ZN(_2300_));
 INV_X1 _6660_ (.A(\aso.z4[6] ),
    .ZN(_2301_));
 AOI21_X1 _6661_ (.A(_2300_),
    .B1(_2301_),
    .B2(\aso.z0[6] ),
    .ZN(_2302_));
 AOI21_X1 _6662_ (.A(_2302_),
    .B1(\aso.z4[7] ),
    .B2(_2273_),
    .ZN(_2303_));
 OR2_X1 _6663_ (.A1(_2281_),
    .A2(_2303_),
    .ZN(_2304_));
 XNOR2_X1 _6664_ (.A(\aso.z0[8] ),
    .B(\aso.z4[8] ),
    .ZN(_2305_));
 XOR2_X1 _6665_ (.A(_2304_),
    .B(_2305_),
    .Z(_2306_));
 NOR2_X1 _6666_ (.A1(_0010_),
    .A2(_2306_),
    .ZN(_2307_));
 NAND2_X1 _6667_ (.A1(_2304_),
    .A2(_2305_),
    .ZN(_2308_));
 OAI21_X1 _6668_ (.A(_2308_),
    .B1(\aso.z4[8] ),
    .B2(_2272_),
    .ZN(_2309_));
 XOR2_X1 _6669_ (.A(\aso.z0[9] ),
    .B(\aso.z4[9] ),
    .Z(_2310_));
 XNOR2_X1 _6670_ (.A(_2309_),
    .B(_2310_),
    .ZN(_2311_));
 NAND2_X1 _6671_ (.A1(\aso.z0[9] ),
    .A2(_2311_),
    .ZN(_2312_));
 XOR2_X1 _6672_ (.A(_2307_),
    .B(_2312_),
    .Z(_2313_));
 INV_X1 _6673_ (.A(\aso.z4[9] ),
    .ZN(_2314_));
 AOI21_X1 _6674_ (.A(_2309_),
    .B1(_2314_),
    .B2(\aso.z0[9] ),
    .ZN(_2315_));
 AOI21_X1 _6675_ (.A(_2315_),
    .B1(\aso.z4[9] ),
    .B2(_2271_),
    .ZN(_2316_));
 XOR2_X1 _6676_ (.A(\aso.z0[10] ),
    .B(\aso.z4[10] ),
    .Z(_2317_));
 XNOR2_X1 _6677_ (.A(_2316_),
    .B(_2317_),
    .ZN(_2318_));
 NAND3_X1 _6678_ (.A1(\aso.z0[4] ),
    .A2(\aso.z0[0] ),
    .A3(_2318_),
    .ZN(_2319_));
 NAND2_X1 _6679_ (.A1(\aso.z0[0] ),
    .A2(_2318_),
    .ZN(_2320_));
 NAND2_X1 _6680_ (.A1(\aso.z0[4] ),
    .A2(_2318_),
    .ZN(_2321_));
 XOR2_X1 _6681_ (.A(_2320_),
    .B(_2321_),
    .Z(_2322_));
 NAND3_X1 _6682_ (.A1(\aso.z0[5] ),
    .A2(_2318_),
    .A3(_2322_),
    .ZN(_2323_));
 NAND2_X1 _6683_ (.A1(_2319_),
    .A2(_2323_),
    .ZN(_2324_));
 NAND2_X1 _6684_ (.A1(\aso.z0[8] ),
    .A2(_2311_),
    .ZN(_2325_));
 OAI21_X1 _6685_ (.A(_2318_),
    .B1(\aso.z0[6] ),
    .B2(\aso.z0[7] ),
    .ZN(_2326_));
 NAND3_X1 _6686_ (.A1(\aso.z0[7] ),
    .A2(\aso.z0[6] ),
    .A3(_2318_),
    .ZN(_2327_));
 INV_X1 _6687_ (.A(_2327_),
    .ZN(_2328_));
 NOR2_X1 _6688_ (.A1(_2326_),
    .A2(_2328_),
    .ZN(_2329_));
 XNOR2_X1 _6689_ (.A(_2325_),
    .B(_2329_),
    .ZN(_2330_));
 AND2_X1 _6690_ (.A1(_2324_),
    .A2(_2330_),
    .ZN(_2331_));
 XOR2_X1 _6691_ (.A(_2324_),
    .B(_2330_),
    .Z(_2332_));
 NAND2_X1 _6692_ (.A1(\aso.z0[7] ),
    .A2(_2311_),
    .ZN(_2333_));
 NAND2_X1 _6693_ (.A1(\aso.z0[6] ),
    .A2(_2318_),
    .ZN(_2334_));
 XOR2_X1 _6694_ (.A(_2333_),
    .B(_2334_),
    .Z(_2335_));
 NAND3_X1 _6695_ (.A1(\aso.z0[8] ),
    .A2(_2306_),
    .A3(_2335_),
    .ZN(_2336_));
 OAI21_X1 _6696_ (.A(_2336_),
    .B1(_2334_),
    .B2(_2333_),
    .ZN(_2337_));
 AOI21_X1 _6697_ (.A(_2331_),
    .B1(_2332_),
    .B2(_2337_),
    .ZN(_2338_));
 NOR2_X1 _6698_ (.A1(_2313_),
    .A2(_2338_),
    .ZN(_2339_));
 XOR2_X1 _6699_ (.A(_2313_),
    .B(_2338_),
    .Z(_2340_));
 XNOR2_X1 _6700_ (.A(\aso.z0[7] ),
    .B(\aso.z4[7] ),
    .ZN(_2341_));
 XNOR2_X1 _6701_ (.A(_2302_),
    .B(_2341_),
    .ZN(_2342_));
 NAND2_X1 _6702_ (.A1(\aso.z0[9] ),
    .A2(_2306_),
    .ZN(_2343_));
 NOR3_X1 _6703_ (.A1(_0010_),
    .A2(_2342_),
    .A3(_2343_),
    .ZN(_2344_));
 AOI21_X1 _6704_ (.A(_2339_),
    .B1(_2340_),
    .B2(_2344_),
    .ZN(_2345_));
 AND3_X1 _6705_ (.A1(\aso.z0[3] ),
    .A2(\aso.z0[2] ),
    .A3(_2318_),
    .ZN(_2346_));
 NAND2_X1 _6706_ (.A1(\aso.z0[1] ),
    .A2(_2346_),
    .ZN(_2347_));
 NAND2_X1 _6707_ (.A1(\aso.z0[5] ),
    .A2(_2318_),
    .ZN(_2348_));
 XOR2_X1 _6708_ (.A(_2322_),
    .B(_2348_),
    .Z(_2349_));
 OR2_X1 _6709_ (.A1(_2347_),
    .A2(_2349_),
    .ZN(_2350_));
 NAND2_X1 _6710_ (.A1(\aso.z0[1] ),
    .A2(_2318_),
    .ZN(_2351_));
 OAI21_X1 _6711_ (.A(_2318_),
    .B1(\aso.z0[2] ),
    .B2(\aso.z0[3] ),
    .ZN(_2352_));
 NAND3_X1 _6712_ (.A1(_2351_),
    .A2(_2352_),
    .A3(_2349_),
    .ZN(_2353_));
 NAND2_X1 _6713_ (.A1(_2350_),
    .A2(_2353_),
    .ZN(_2354_));
 XNOR2_X1 _6714_ (.A(_2337_),
    .B(_2332_),
    .ZN(_2355_));
 OAI21_X1 _6715_ (.A(_2350_),
    .B1(_2354_),
    .B2(_2355_),
    .ZN(_2356_));
 NAND2_X1 _6716_ (.A1(\aso.z0[8] ),
    .A2(_2318_),
    .ZN(_2357_));
 XOR2_X1 _6717_ (.A(_2329_),
    .B(_2357_),
    .Z(_2358_));
 XOR2_X1 _6718_ (.A(_2324_),
    .B(_2358_),
    .Z(_2359_));
 NAND3_X1 _6719_ (.A1(\aso.z0[8] ),
    .A2(_2311_),
    .A3(_2329_),
    .ZN(_2360_));
 AOI21_X1 _6720_ (.A(_2359_),
    .B1(_2360_),
    .B2(_2327_),
    .ZN(_2361_));
 AND3_X1 _6721_ (.A1(_2327_),
    .A2(_2360_),
    .A3(_2359_),
    .ZN(_2362_));
 OR2_X1 _6722_ (.A1(_2361_),
    .A2(_2362_),
    .ZN(_2363_));
 XNOR2_X1 _6723_ (.A(_2354_),
    .B(_2363_),
    .ZN(_2364_));
 INV_X1 _6724_ (.A(_2364_),
    .ZN(_2365_));
 NAND2_X1 _6725_ (.A1(_2356_),
    .A2(_2365_),
    .ZN(_2366_));
 XOR2_X1 _6726_ (.A(_2356_),
    .B(_2364_),
    .Z(_2367_));
 XNOR2_X1 _6727_ (.A(_2344_),
    .B(_2340_),
    .ZN(_2368_));
 OAI21_X1 _6728_ (.A(_2366_),
    .B1(_2367_),
    .B2(_2368_),
    .ZN(_2369_));
 NAND3_X1 _6729_ (.A1(\aso.z0[9] ),
    .A2(_2311_),
    .A3(_2307_),
    .ZN(_2370_));
 NOR2_X1 _6730_ (.A1(_0010_),
    .A2(_2311_),
    .ZN(_2371_));
 NAND2_X1 _6731_ (.A1(\aso.z0[9] ),
    .A2(_2318_),
    .ZN(_2372_));
 XOR2_X1 _6732_ (.A(_2371_),
    .B(_2372_),
    .Z(_2373_));
 AOI21_X1 _6733_ (.A(_2358_),
    .B1(_2323_),
    .B2(_2319_),
    .ZN(_2374_));
 NOR2_X1 _6734_ (.A1(_2374_),
    .A2(_2361_),
    .ZN(_2375_));
 XNOR2_X1 _6735_ (.A(_2373_),
    .B(_2375_),
    .ZN(_2376_));
 XOR2_X1 _6736_ (.A(_2370_),
    .B(_2376_),
    .Z(_2377_));
 NAND3_X1 _6737_ (.A1(\aso.z0[8] ),
    .A2(_2318_),
    .A3(_2329_),
    .ZN(_2378_));
 AOI21_X1 _6738_ (.A(_2359_),
    .B1(_2378_),
    .B2(_2327_),
    .ZN(_2379_));
 AND3_X1 _6739_ (.A1(_2327_),
    .A2(_2378_),
    .A3(_2359_),
    .ZN(_2380_));
 OR2_X1 _6740_ (.A1(_2379_),
    .A2(_2380_),
    .ZN(_2381_));
 XNOR2_X1 _6741_ (.A(_2354_),
    .B(_2381_),
    .ZN(_2382_));
 OR2_X1 _6742_ (.A1(_2354_),
    .A2(_2363_),
    .ZN(_2383_));
 AOI21_X1 _6743_ (.A(_2382_),
    .B1(_2383_),
    .B2(_2350_),
    .ZN(_2384_));
 AND3_X1 _6744_ (.A1(_2350_),
    .A2(_2383_),
    .A3(_2382_),
    .ZN(_2385_));
 NOR2_X1 _6745_ (.A1(_2384_),
    .A2(_2385_),
    .ZN(_2386_));
 XNOR2_X1 _6746_ (.A(_2377_),
    .B(_2386_),
    .ZN(_2387_));
 XNOR2_X1 _6747_ (.A(_2369_),
    .B(_2387_),
    .ZN(_2388_));
 XOR2_X1 _6748_ (.A(_2345_),
    .B(_2388_),
    .Z(_2389_));
 NOR2_X1 _6749_ (.A1(_0010_),
    .A2(_2342_),
    .ZN(_2390_));
 XOR2_X1 _6750_ (.A(_2390_),
    .B(_2343_),
    .Z(_2391_));
 NAND2_X1 _6751_ (.A1(\aso.z0[8] ),
    .A2(_2306_),
    .ZN(_2392_));
 XNOR2_X1 _6752_ (.A(_2392_),
    .B(_2335_),
    .ZN(_2393_));
 AND2_X1 _6753_ (.A1(_2393_),
    .A2(_2324_),
    .ZN(_2394_));
 XOR2_X1 _6754_ (.A(_2393_),
    .B(_2324_),
    .Z(_2395_));
 NAND2_X1 _6755_ (.A1(\aso.z0[7] ),
    .A2(_2306_),
    .ZN(_2396_));
 NAND2_X1 _6756_ (.A1(\aso.z0[6] ),
    .A2(_2311_),
    .ZN(_2397_));
 XOR2_X1 _6757_ (.A(_2396_),
    .B(_2397_),
    .Z(_2398_));
 NAND3_X1 _6758_ (.A1(\aso.z0[8] ),
    .A2(_2342_),
    .A3(_2398_),
    .ZN(_2399_));
 OAI21_X1 _6759_ (.A(_2399_),
    .B1(_2397_),
    .B2(_2396_),
    .ZN(_2400_));
 AOI21_X1 _6760_ (.A(_2394_),
    .B1(_2395_),
    .B2(_2400_),
    .ZN(_2401_));
 OR2_X1 _6761_ (.A1(_2391_),
    .A2(_2401_),
    .ZN(_2402_));
 XNOR2_X1 _6762_ (.A(_2391_),
    .B(_2401_),
    .ZN(_2403_));
 XOR2_X1 _6763_ (.A(_2282_),
    .B(_2299_),
    .Z(_2404_));
 NAND2_X1 _6764_ (.A1(\aso.z0[9] ),
    .A2(_2342_),
    .ZN(_2405_));
 OR3_X1 _6765_ (.A1(_0010_),
    .A2(_2404_),
    .A3(_2405_),
    .ZN(_2406_));
 OAI21_X1 _6766_ (.A(_2402_),
    .B1(_2403_),
    .B2(_2406_),
    .ZN(_2407_));
 XNOR2_X1 _6767_ (.A(_2400_),
    .B(_2395_),
    .ZN(_2408_));
 OR2_X1 _6768_ (.A1(_2408_),
    .A2(_2354_),
    .ZN(_2409_));
 AND2_X1 _6769_ (.A1(_2350_),
    .A2(_2409_),
    .ZN(_2410_));
 XNOR2_X1 _6770_ (.A(_2354_),
    .B(_2355_),
    .ZN(_2411_));
 NOR2_X1 _6771_ (.A1(_2410_),
    .A2(_2411_),
    .ZN(_2412_));
 XNOR2_X1 _6772_ (.A(_2406_),
    .B(_2403_),
    .ZN(_2413_));
 XNOR2_X1 _6773_ (.A(_2410_),
    .B(_2411_),
    .ZN(_2414_));
 NOR2_X1 _6774_ (.A1(_2413_),
    .A2(_2414_),
    .ZN(_2415_));
 NOR2_X1 _6775_ (.A1(_2412_),
    .A2(_2415_),
    .ZN(_2416_));
 XOR2_X1 _6776_ (.A(_2368_),
    .B(_2367_),
    .Z(_2417_));
 XNOR2_X1 _6777_ (.A(_2416_),
    .B(_2417_),
    .ZN(_2418_));
 NAND2_X1 _6778_ (.A1(_2407_),
    .A2(_2418_),
    .ZN(_2419_));
 OAI21_X1 _6779_ (.A(_2417_),
    .B1(_2415_),
    .B2(_2412_),
    .ZN(_2420_));
 AOI21_X1 _6780_ (.A(_2389_),
    .B1(_2419_),
    .B2(_2420_),
    .ZN(_2421_));
 AND3_X1 _6781_ (.A1(_2420_),
    .A2(_2419_),
    .A3(_2389_),
    .ZN(_2422_));
 NOR2_X1 _6782_ (.A1(_2421_),
    .A2(_2422_),
    .ZN(_2423_));
 INV_X1 _6783_ (.A(_2423_),
    .ZN(_2424_));
 NAND2_X1 _6784_ (.A1(_2351_),
    .A2(_2352_),
    .ZN(_2425_));
 NAND2_X1 _6785_ (.A1(_2347_),
    .A2(_2425_),
    .ZN(_2426_));
 XOR2_X1 _6786_ (.A(_2349_),
    .B(_2426_),
    .Z(_2427_));
 NAND2_X1 _6787_ (.A1(\aso.z0[5] ),
    .A2(_2311_),
    .ZN(_2428_));
 XOR2_X1 _6788_ (.A(_2322_),
    .B(_2428_),
    .Z(_2429_));
 OAI21_X1 _6789_ (.A(_2347_),
    .B1(_2426_),
    .B2(_2429_),
    .ZN(_2430_));
 NAND2_X1 _6790_ (.A1(_2427_),
    .A2(_2430_),
    .ZN(_2431_));
 NAND2_X1 _6791_ (.A1(\aso.z0[8] ),
    .A2(_2342_),
    .ZN(_2432_));
 XNOR2_X1 _6792_ (.A(_2432_),
    .B(_2398_),
    .ZN(_2433_));
 NAND3_X1 _6793_ (.A1(\aso.z0[5] ),
    .A2(_2322_),
    .A3(_2311_),
    .ZN(_2434_));
 NAND2_X1 _6794_ (.A1(_2319_),
    .A2(_2434_),
    .ZN(_2435_));
 XOR2_X1 _6795_ (.A(_2433_),
    .B(_2435_),
    .Z(_2436_));
 INV_X1 _6796_ (.A(_2404_),
    .ZN(_2437_));
 NAND2_X1 _6797_ (.A1(\aso.z0[6] ),
    .A2(_2342_),
    .ZN(_2438_));
 NOR2_X1 _6798_ (.A1(_2396_),
    .A2(_2438_),
    .ZN(_2439_));
 AOI22_X1 _6799_ (.A1(\aso.z0[6] ),
    .A2(_2306_),
    .B1(_2342_),
    .B2(\aso.z0[7] ),
    .ZN(_2440_));
 NOR4_X1 _6800_ (.A1(_2272_),
    .A2(_2437_),
    .A3(_2439_),
    .A4(_2440_),
    .ZN(_2441_));
 OAI21_X1 _6801_ (.A(_2436_),
    .B1(_2441_),
    .B2(_2439_),
    .ZN(_2442_));
 OR3_X1 _6802_ (.A1(_2439_),
    .A2(_2441_),
    .A3(_2436_),
    .ZN(_2443_));
 NAND2_X1 _6803_ (.A1(_2442_),
    .A2(_2443_),
    .ZN(_2444_));
 NOR2_X1 _6804_ (.A1(_2427_),
    .A2(_2430_),
    .ZN(_2445_));
 OAI21_X1 _6805_ (.A(_2431_),
    .B1(_2444_),
    .B2(_2445_),
    .ZN(_2446_));
 XOR2_X1 _6806_ (.A(_2408_),
    .B(_2354_),
    .Z(_2447_));
 NAND2_X1 _6807_ (.A1(_2446_),
    .A2(_2447_),
    .ZN(_2448_));
 XOR2_X1 _6808_ (.A(_2283_),
    .B(_2296_),
    .Z(_2449_));
 OR4_X1 _6809_ (.A1(_2271_),
    .A2(_0010_),
    .A3(_2437_),
    .A4(_2449_),
    .ZN(_2450_));
 OAI21_X1 _6810_ (.A(_2405_),
    .B1(_2404_),
    .B2(_0010_),
    .ZN(_2451_));
 NAND2_X1 _6811_ (.A1(_2406_),
    .A2(_2451_),
    .ZN(_2452_));
 NAND2_X1 _6812_ (.A1(_2433_),
    .A2(_2435_),
    .ZN(_2453_));
 NAND2_X1 _6813_ (.A1(_2453_),
    .A2(_2442_),
    .ZN(_2454_));
 XOR2_X1 _6814_ (.A(_2452_),
    .B(_2454_),
    .Z(_2455_));
 XNOR2_X1 _6815_ (.A(_2450_),
    .B(_2455_),
    .ZN(_2456_));
 XNOR2_X1 _6816_ (.A(_2446_),
    .B(_2447_),
    .ZN(_2457_));
 OAI21_X1 _6817_ (.A(_2448_),
    .B1(_2456_),
    .B2(_2457_),
    .ZN(_2458_));
 XNOR2_X1 _6818_ (.A(_2413_),
    .B(_2414_),
    .ZN(_2459_));
 INV_X1 _6819_ (.A(_2459_),
    .ZN(_2460_));
 NAND2_X1 _6820_ (.A1(_2458_),
    .A2(_2460_),
    .ZN(_2461_));
 NAND3_X1 _6821_ (.A1(_2406_),
    .A2(_2451_),
    .A3(_2454_),
    .ZN(_2462_));
 OAI21_X1 _6822_ (.A(_2462_),
    .B1(_2455_),
    .B2(_2450_),
    .ZN(_2463_));
 INV_X1 _6823_ (.A(_2463_),
    .ZN(_2464_));
 XOR2_X1 _6824_ (.A(_2458_),
    .B(_2459_),
    .Z(_2465_));
 OAI21_X1 _6825_ (.A(_2461_),
    .B1(_2464_),
    .B2(_2465_),
    .ZN(_2466_));
 XNOR2_X1 _6826_ (.A(_2407_),
    .B(_2418_),
    .ZN(_2467_));
 INV_X1 _6827_ (.A(_2467_),
    .ZN(_2468_));
 NAND2_X1 _6828_ (.A1(_2466_),
    .A2(_2468_),
    .ZN(_2469_));
 XNOR2_X1 _6829_ (.A(_2464_),
    .B(_2465_),
    .ZN(_2470_));
 OAI22_X1 _6830_ (.A1(_2271_),
    .A2(_2437_),
    .B1(_2449_),
    .B2(_0010_),
    .ZN(_2471_));
 NAND2_X1 _6831_ (.A1(_2450_),
    .A2(_2471_),
    .ZN(_2472_));
 NAND2_X1 _6832_ (.A1(\aso.z0[7] ),
    .A2(_2404_),
    .ZN(_2473_));
 XOR2_X1 _6833_ (.A(_2438_),
    .B(_2473_),
    .Z(_2474_));
 NAND3_X1 _6834_ (.A1(\aso.z0[8] ),
    .A2(_2449_),
    .A3(_2474_),
    .ZN(_2475_));
 OAI21_X1 _6835_ (.A(_2475_),
    .B1(_2473_),
    .B2(_2438_),
    .ZN(_2476_));
 NOR2_X1 _6836_ (.A1(_2439_),
    .A2(_2440_),
    .ZN(_2477_));
 AOI21_X1 _6837_ (.A(_2477_),
    .B1(_2404_),
    .B2(\aso.z0[8] ),
    .ZN(_2478_));
 NOR2_X1 _6838_ (.A1(_2441_),
    .A2(_2478_),
    .ZN(_2479_));
 NAND2_X1 _6839_ (.A1(\aso.z0[0] ),
    .A2(_2311_),
    .ZN(_2480_));
 NAND2_X1 _6840_ (.A1(\aso.z0[4] ),
    .A2(_2311_),
    .ZN(_2481_));
 XNOR2_X1 _6841_ (.A(_2320_),
    .B(_2481_),
    .ZN(_2482_));
 NAND2_X1 _6842_ (.A1(\aso.z0[5] ),
    .A2(_2306_),
    .ZN(_2483_));
 OAI22_X1 _6843_ (.A1(_2321_),
    .A2(_2480_),
    .B1(_2482_),
    .B2(_2483_),
    .ZN(_2484_));
 XOR2_X1 _6844_ (.A(_2479_),
    .B(_2484_),
    .Z(_2485_));
 NAND2_X1 _6845_ (.A1(_2476_),
    .A2(_2485_),
    .ZN(_2486_));
 NAND2_X1 _6846_ (.A1(_2479_),
    .A2(_2484_),
    .ZN(_2487_));
 AOI21_X1 _6847_ (.A(_2472_),
    .B1(_2486_),
    .B2(_2487_),
    .ZN(_2488_));
 INV_X1 _6848_ (.A(_2488_),
    .ZN(_2489_));
 NAND3_X1 _6849_ (.A1(_2487_),
    .A2(_2486_),
    .A3(_2472_),
    .ZN(_2490_));
 NAND2_X1 _6850_ (.A1(_2489_),
    .A2(_2490_),
    .ZN(_2491_));
 XOR2_X1 _6851_ (.A(_2294_),
    .B(_2295_),
    .Z(_2492_));
 NAND2_X1 _6852_ (.A1(\aso.z0[9] ),
    .A2(_2449_),
    .ZN(_2493_));
 OR3_X1 _6853_ (.A1(_0010_),
    .A2(_2492_),
    .A3(_2493_),
    .ZN(_2494_));
 OAI21_X1 _6854_ (.A(_2489_),
    .B1(_2491_),
    .B2(_2494_),
    .ZN(_2495_));
 XOR2_X1 _6855_ (.A(_2427_),
    .B(_2430_),
    .Z(_2496_));
 XNOR2_X1 _6856_ (.A(_2444_),
    .B(_2496_),
    .ZN(_2497_));
 XNOR2_X1 _6857_ (.A(_2476_),
    .B(_2485_),
    .ZN(_2498_));
 NOR2_X1 _6858_ (.A1(_2346_),
    .A2(_2352_),
    .ZN(_2499_));
 XNOR2_X1 _6859_ (.A(_2351_),
    .B(_2499_),
    .ZN(_2500_));
 INV_X1 _6860_ (.A(_0011_),
    .ZN(_2501_));
 AND4_X1 _6861_ (.A1(\aso.z0[2] ),
    .A2(_2501_),
    .A3(_2318_),
    .A4(_2311_),
    .ZN(_2502_));
 AOI22_X1 _6862_ (.A1(\aso.z0[2] ),
    .A2(_2318_),
    .B1(_2311_),
    .B2(_2501_),
    .ZN(_2503_));
 NOR3_X1 _6863_ (.A1(_2351_),
    .A2(_2502_),
    .A3(_2503_),
    .ZN(_2504_));
 OR2_X1 _6864_ (.A1(_2502_),
    .A2(_2504_),
    .ZN(_2505_));
 AND2_X1 _6865_ (.A1(_2500_),
    .A2(_2505_),
    .ZN(_2506_));
 XOR2_X1 _6866_ (.A(_2483_),
    .B(_2482_),
    .Z(_2507_));
 XOR2_X1 _6867_ (.A(_2500_),
    .B(_2505_),
    .Z(_2508_));
 AOI21_X1 _6868_ (.A(_2506_),
    .B1(_2507_),
    .B2(_2508_),
    .ZN(_2509_));
 XOR2_X1 _6869_ (.A(_2426_),
    .B(_2429_),
    .Z(_2510_));
 INV_X1 _6870_ (.A(_2510_),
    .ZN(_2511_));
 XNOR2_X1 _6871_ (.A(_2509_),
    .B(_2511_),
    .ZN(_2512_));
 NOR2_X1 _6872_ (.A1(_2498_),
    .A2(_2512_),
    .ZN(_2513_));
 NOR2_X1 _6873_ (.A1(_2509_),
    .A2(_2511_),
    .ZN(_2514_));
 OAI21_X1 _6874_ (.A(_2497_),
    .B1(_2513_),
    .B2(_2514_),
    .ZN(_2515_));
 XNOR2_X1 _6875_ (.A(_2494_),
    .B(_2491_),
    .ZN(_2516_));
 OR3_X1 _6876_ (.A1(_2514_),
    .A2(_2513_),
    .A3(_2497_),
    .ZN(_2517_));
 NAND2_X1 _6877_ (.A1(_2515_),
    .A2(_2517_),
    .ZN(_2518_));
 OAI21_X1 _6878_ (.A(_2515_),
    .B1(_2516_),
    .B2(_2518_),
    .ZN(_2519_));
 XOR2_X1 _6879_ (.A(_2456_),
    .B(_2457_),
    .Z(_2520_));
 XNOR2_X1 _6880_ (.A(_2519_),
    .B(_2520_),
    .ZN(_2521_));
 INV_X1 _6881_ (.A(_2521_),
    .ZN(_2522_));
 NAND2_X1 _6882_ (.A1(_2495_),
    .A2(_2522_),
    .ZN(_2523_));
 NAND2_X1 _6883_ (.A1(_2519_),
    .A2(_2520_),
    .ZN(_2524_));
 AOI21_X1 _6884_ (.A(_2470_),
    .B1(_2523_),
    .B2(_2524_),
    .ZN(_2525_));
 AND3_X1 _6885_ (.A1(_2524_),
    .A2(_2523_),
    .A3(_2470_),
    .ZN(_2526_));
 NOR2_X1 _6886_ (.A1(_2525_),
    .A2(_2526_),
    .ZN(_2527_));
 XOR2_X1 _6887_ (.A(_2498_),
    .B(_2512_),
    .Z(_2528_));
 NAND2_X1 _6888_ (.A1(\aso.z0[6] ),
    .A2(_2449_),
    .ZN(_2529_));
 NAND2_X1 _6889_ (.A1(\aso.z0[8] ),
    .A2(_2492_),
    .ZN(_2530_));
 INV_X1 _6890_ (.A(_2449_),
    .ZN(_2531_));
 OAI22_X1 _6891_ (.A1(_2274_),
    .A2(_2437_),
    .B1(_2531_),
    .B2(_2273_),
    .ZN(_2532_));
 OAI21_X1 _6892_ (.A(_2532_),
    .B1(_2529_),
    .B2(_2473_),
    .ZN(_2533_));
 OAI22_X1 _6893_ (.A1(_2473_),
    .A2(_2529_),
    .B1(_2530_),
    .B2(_2533_),
    .ZN(_2534_));
 NAND2_X1 _6894_ (.A1(\aso.z0[8] ),
    .A2(_2449_),
    .ZN(_2535_));
 XNOR2_X1 _6895_ (.A(_2535_),
    .B(_2474_),
    .ZN(_2536_));
 NAND2_X1 _6896_ (.A1(\aso.z0[4] ),
    .A2(_2306_),
    .ZN(_2537_));
 XOR2_X1 _6897_ (.A(_2320_),
    .B(_2537_),
    .Z(_2538_));
 NAND3_X1 _6898_ (.A1(\aso.z0[5] ),
    .A2(_2342_),
    .A3(_2538_),
    .ZN(_2539_));
 OAI21_X1 _6899_ (.A(_2539_),
    .B1(_2537_),
    .B2(_2320_),
    .ZN(_2540_));
 XOR2_X1 _6900_ (.A(_2536_),
    .B(_2540_),
    .Z(_2541_));
 XNOR2_X1 _6901_ (.A(_2534_),
    .B(_2541_),
    .ZN(_2542_));
 XNOR2_X1 _6902_ (.A(_2507_),
    .B(_2508_),
    .ZN(_2543_));
 NAND2_X1 _6903_ (.A1(\aso.z0[5] ),
    .A2(_2342_),
    .ZN(_2544_));
 XNOR2_X1 _6904_ (.A(_2544_),
    .B(_2538_),
    .ZN(_2545_));
 AND4_X1 _6905_ (.A1(\aso.z0[3] ),
    .A2(\aso.z0[2] ),
    .A3(_2306_),
    .A4(_2311_),
    .ZN(_2546_));
 AOI22_X1 _6906_ (.A1(\aso.z0[3] ),
    .A2(_2306_),
    .B1(_2311_),
    .B2(\aso.z0[2] ),
    .ZN(_2547_));
 OR2_X1 _6907_ (.A1(_2546_),
    .A2(_2547_),
    .ZN(_2548_));
 NOR2_X1 _6908_ (.A1(_2351_),
    .A2(_2548_),
    .ZN(_2549_));
 OR2_X1 _6909_ (.A1(_2546_),
    .A2(_2549_),
    .ZN(_2550_));
 OR3_X1 _6910_ (.A1(_2351_),
    .A2(_2502_),
    .A3(_2503_),
    .ZN(_2551_));
 OAI21_X1 _6911_ (.A(_2351_),
    .B1(_2502_),
    .B2(_2503_),
    .ZN(_2552_));
 AND2_X1 _6912_ (.A1(_2551_),
    .A2(_2552_),
    .ZN(_2553_));
 XNOR2_X1 _6913_ (.A(_2550_),
    .B(_2553_),
    .ZN(_2554_));
 INV_X1 _6914_ (.A(_2554_),
    .ZN(_2555_));
 NAND2_X1 _6915_ (.A1(_2545_),
    .A2(_2555_),
    .ZN(_2556_));
 NAND2_X1 _6916_ (.A1(_2550_),
    .A2(_2553_),
    .ZN(_2557_));
 AOI21_X1 _6917_ (.A(_2543_),
    .B1(_2556_),
    .B2(_2557_),
    .ZN(_2558_));
 AND3_X1 _6918_ (.A1(_2557_),
    .A2(_2556_),
    .A3(_2543_),
    .ZN(_2559_));
 OR2_X1 _6919_ (.A1(_2558_),
    .A2(_2559_),
    .ZN(_2560_));
 NOR2_X1 _6920_ (.A1(_2542_),
    .A2(_2560_),
    .ZN(_2561_));
 OAI21_X1 _6921_ (.A(_2528_),
    .B1(_2561_),
    .B2(_2558_),
    .ZN(_2562_));
 OR3_X1 _6922_ (.A1(_2558_),
    .A2(_2561_),
    .A3(_2528_),
    .ZN(_2563_));
 NAND2_X1 _6923_ (.A1(_2562_),
    .A2(_2563_),
    .ZN(_2564_));
 INV_X1 _6924_ (.A(_2492_),
    .ZN(_2565_));
 XOR2_X1 _6925_ (.A(_2286_),
    .B(_2293_),
    .Z(_2566_));
 OR4_X1 _6926_ (.A1(_2271_),
    .A2(_0010_),
    .A3(_2565_),
    .A4(_2566_),
    .ZN(_2567_));
 OAI21_X1 _6927_ (.A(_2493_),
    .B1(_2492_),
    .B2(_0010_),
    .ZN(_2568_));
 NAND2_X1 _6928_ (.A1(_2494_),
    .A2(_2568_),
    .ZN(_2569_));
 AOI22_X1 _6929_ (.A1(_2536_),
    .A2(_2540_),
    .B1(_2541_),
    .B2(_2534_),
    .ZN(_2570_));
 XNOR2_X1 _6930_ (.A(_2569_),
    .B(_2570_),
    .ZN(_2571_));
 XNOR2_X1 _6931_ (.A(_2567_),
    .B(_2571_),
    .ZN(_2572_));
 OAI21_X1 _6932_ (.A(_2562_),
    .B1(_2564_),
    .B2(_2572_),
    .ZN(_2573_));
 XNOR2_X1 _6933_ (.A(_2516_),
    .B(_2518_),
    .ZN(_2574_));
 INV_X1 _6934_ (.A(_2574_),
    .ZN(_2575_));
 NAND2_X1 _6935_ (.A1(_2573_),
    .A2(_2575_),
    .ZN(_2576_));
 XNOR2_X1 _6936_ (.A(_2573_),
    .B(_2575_),
    .ZN(_2577_));
 OR2_X1 _6937_ (.A1(_2567_),
    .A2(_2571_),
    .ZN(_2578_));
 OAI21_X1 _6938_ (.A(_2578_),
    .B1(_2570_),
    .B2(_2569_),
    .ZN(_2579_));
 INV_X1 _6939_ (.A(_2579_),
    .ZN(_2580_));
 OAI21_X1 _6940_ (.A(_2576_),
    .B1(_2577_),
    .B2(_2580_),
    .ZN(_2581_));
 INV_X1 _6941_ (.A(_2581_),
    .ZN(_2582_));
 XOR2_X1 _6942_ (.A(_2495_),
    .B(_2521_),
    .Z(_2583_));
 NOR2_X1 _6943_ (.A1(_2582_),
    .A2(_2583_),
    .ZN(_2584_));
 AND2_X1 _6944_ (.A1(_2527_),
    .A2(_2584_),
    .ZN(_2585_));
 AND2_X1 _6945_ (.A1(\aso.z0[3] ),
    .A2(_2342_),
    .ZN(_2586_));
 XNOR2_X1 _6946_ (.A(_0010_),
    .B(_2586_),
    .ZN(_2587_));
 AND3_X1 _6947_ (.A1(\aso.z0[2] ),
    .A2(_2306_),
    .A3(_2587_),
    .ZN(_2588_));
 AOI21_X1 _6948_ (.A(_2588_),
    .B1(_2586_),
    .B2(\aso.z0[10] ),
    .ZN(_2589_));
 INV_X1 _6949_ (.A(_2589_),
    .ZN(_2590_));
 XOR2_X1 _6950_ (.A(_2351_),
    .B(_2548_),
    .Z(_2591_));
 NAND2_X1 _6951_ (.A1(\aso.z0[5] ),
    .A2(_2404_),
    .ZN(_2592_));
 NAND2_X1 _6952_ (.A1(\aso.z0[4] ),
    .A2(_2342_),
    .ZN(_2593_));
 XNOR2_X1 _6953_ (.A(_2320_),
    .B(_2593_),
    .ZN(_2594_));
 XOR2_X1 _6954_ (.A(_2592_),
    .B(_2594_),
    .Z(_2595_));
 XNOR2_X1 _6955_ (.A(_2589_),
    .B(_2591_),
    .ZN(_2596_));
 AOI22_X1 _6956_ (.A1(_2590_),
    .A2(_2591_),
    .B1(_2595_),
    .B2(_2596_),
    .ZN(_2597_));
 XOR2_X1 _6957_ (.A(_2545_),
    .B(_2554_),
    .Z(_2598_));
 OR2_X1 _6958_ (.A1(_2597_),
    .A2(_2598_),
    .ZN(_2599_));
 NAND2_X1 _6959_ (.A1(\aso.z0[7] ),
    .A2(_2492_),
    .ZN(_2600_));
 XOR2_X1 _6960_ (.A(_2529_),
    .B(_2600_),
    .Z(_2601_));
 NAND3_X1 _6961_ (.A1(\aso.z0[8] ),
    .A2(_2566_),
    .A3(_2601_),
    .ZN(_2602_));
 OAI21_X1 _6962_ (.A(_2602_),
    .B1(_2600_),
    .B2(_2529_),
    .ZN(_2603_));
 XOR2_X1 _6963_ (.A(_2530_),
    .B(_2533_),
    .Z(_2604_));
 NAND2_X1 _6964_ (.A1(\aso.z0[0] ),
    .A2(_2342_),
    .ZN(_2605_));
 OAI22_X1 _6965_ (.A1(_2321_),
    .A2(_2605_),
    .B1(_2594_),
    .B2(_2592_),
    .ZN(_2606_));
 XOR2_X1 _6966_ (.A(_2604_),
    .B(_2606_),
    .Z(_2607_));
 XNOR2_X1 _6967_ (.A(_2603_),
    .B(_2607_),
    .ZN(_2608_));
 AND2_X1 _6968_ (.A1(_2597_),
    .A2(_2598_),
    .ZN(_2609_));
 OAI21_X1 _6969_ (.A(_2599_),
    .B1(_2608_),
    .B2(_2609_),
    .ZN(_2610_));
 XOR2_X1 _6970_ (.A(_2542_),
    .B(_2560_),
    .Z(_2611_));
 NAND2_X1 _6971_ (.A1(_2610_),
    .A2(_2611_),
    .ZN(_2612_));
 INV_X1 _6972_ (.A(_2566_),
    .ZN(_2613_));
 XOR2_X1 _6973_ (.A(_2291_),
    .B(_2292_),
    .Z(_2614_));
 OR4_X1 _6974_ (.A1(_2271_),
    .A2(_0010_),
    .A3(_2613_),
    .A4(_2614_),
    .ZN(_2615_));
 OAI22_X1 _6975_ (.A1(_2271_),
    .A2(_2565_),
    .B1(_2566_),
    .B2(_0010_),
    .ZN(_2616_));
 NAND2_X1 _6976_ (.A1(_2567_),
    .A2(_2616_),
    .ZN(_2617_));
 NAND2_X1 _6977_ (.A1(_2603_),
    .A2(_2607_),
    .ZN(_2618_));
 NAND2_X1 _6978_ (.A1(_2604_),
    .A2(_2606_),
    .ZN(_2619_));
 AOI21_X1 _6979_ (.A(_2617_),
    .B1(_2618_),
    .B2(_2619_),
    .ZN(_2620_));
 AND3_X1 _6980_ (.A1(_2619_),
    .A2(_2618_),
    .A3(_2617_),
    .ZN(_2621_));
 OR2_X1 _6981_ (.A1(_2620_),
    .A2(_2621_),
    .ZN(_2622_));
 XOR2_X1 _6982_ (.A(_2615_),
    .B(_2622_),
    .Z(_2623_));
 INV_X1 _6983_ (.A(_2623_),
    .ZN(_2624_));
 XNOR2_X1 _6984_ (.A(_2610_),
    .B(_2611_),
    .ZN(_2625_));
 OAI21_X1 _6985_ (.A(_2612_),
    .B1(_2624_),
    .B2(_2625_),
    .ZN(_2626_));
 XOR2_X1 _6986_ (.A(_2572_),
    .B(_2564_),
    .Z(_2627_));
 NAND2_X1 _6987_ (.A1(_2626_),
    .A2(_2627_),
    .ZN(_2628_));
 INV_X1 _6988_ (.A(_2620_),
    .ZN(_2629_));
 OAI21_X1 _6989_ (.A(_2629_),
    .B1(_2621_),
    .B2(_2615_),
    .ZN(_2630_));
 INV_X1 _6990_ (.A(_2630_),
    .ZN(_2631_));
 XNOR2_X1 _6991_ (.A(_2626_),
    .B(_2627_),
    .ZN(_2632_));
 OAI21_X1 _6992_ (.A(_2628_),
    .B1(_2631_),
    .B2(_2632_),
    .ZN(_2633_));
 XNOR2_X1 _6993_ (.A(_2580_),
    .B(_2577_),
    .ZN(_2634_));
 XOR2_X1 _6994_ (.A(_2633_),
    .B(_2634_),
    .Z(_2635_));
 XNOR2_X1 _6995_ (.A(_2624_),
    .B(_2625_),
    .ZN(_2636_));
 XOR2_X1 _6996_ (.A(_2288_),
    .B(_2289_),
    .Z(_2637_));
 NAND2_X1 _6997_ (.A1(\aso.z0[9] ),
    .A2(_2614_),
    .ZN(_2638_));
 OR3_X1 _6998_ (.A1(_0010_),
    .A2(_2637_),
    .A3(_2638_),
    .ZN(_2639_));
 OAI22_X1 _6999_ (.A1(_2271_),
    .A2(_2613_),
    .B1(_2614_),
    .B2(_0010_),
    .ZN(_2640_));
 NAND2_X1 _7000_ (.A1(_2615_),
    .A2(_2640_),
    .ZN(_2641_));
 NAND2_X1 _7001_ (.A1(\aso.z0[8] ),
    .A2(_2566_),
    .ZN(_2642_));
 XNOR2_X1 _7002_ (.A(_2642_),
    .B(_2601_),
    .ZN(_2643_));
 NAND2_X1 _7003_ (.A1(\aso.z0[1] ),
    .A2(_2311_),
    .ZN(_2644_));
 XOR2_X1 _7004_ (.A(_2320_),
    .B(_2644_),
    .Z(_2645_));
 NAND3_X1 _7005_ (.A1(\aso.z0[4] ),
    .A2(_2404_),
    .A3(_2645_),
    .ZN(_2646_));
 OAI21_X1 _7006_ (.A(_2646_),
    .B1(_2480_),
    .B2(_2351_),
    .ZN(_2647_));
 AND2_X1 _7007_ (.A1(_2643_),
    .A2(_2647_),
    .ZN(_2648_));
 XOR2_X1 _7008_ (.A(_2643_),
    .B(_2647_),
    .Z(_2649_));
 NAND2_X1 _7009_ (.A1(\aso.z0[5] ),
    .A2(_2492_),
    .ZN(_2650_));
 NAND2_X1 _7010_ (.A1(\aso.z0[7] ),
    .A2(_2566_),
    .ZN(_2651_));
 AOI22_X1 _7011_ (.A1(\aso.z0[5] ),
    .A2(_2449_),
    .B1(_2492_),
    .B2(\aso.z0[6] ),
    .ZN(_2652_));
 OAI22_X1 _7012_ (.A1(_2529_),
    .A2(_2650_),
    .B1(_2651_),
    .B2(_2652_),
    .ZN(_2653_));
 AOI21_X1 _7013_ (.A(_2648_),
    .B1(_2649_),
    .B2(_2653_),
    .ZN(_2654_));
 XNOR2_X1 _7014_ (.A(_2641_),
    .B(_2654_),
    .ZN(_2655_));
 XOR2_X1 _7015_ (.A(_2639_),
    .B(_2655_),
    .Z(_2656_));
 XOR2_X1 _7016_ (.A(_2597_),
    .B(_2598_),
    .Z(_2657_));
 XNOR2_X1 _7017_ (.A(_2608_),
    .B(_2657_),
    .ZN(_2658_));
 XNOR2_X1 _7018_ (.A(_2653_),
    .B(_2649_),
    .ZN(_2659_));
 NAND2_X1 _7019_ (.A1(\aso.z0[4] ),
    .A2(_2404_),
    .ZN(_2660_));
 XOR2_X1 _7020_ (.A(_2660_),
    .B(_2645_),
    .Z(_2661_));
 NAND4_X1 _7021_ (.A1(\aso.z0[2] ),
    .A2(_2501_),
    .A3(_2342_),
    .A4(_2404_),
    .ZN(_2662_));
 NAND2_X1 _7022_ (.A1(\aso.z0[2] ),
    .A2(_2342_),
    .ZN(_2663_));
 OAI21_X1 _7023_ (.A(_2663_),
    .B1(_2437_),
    .B2(_0011_),
    .ZN(_2664_));
 NAND2_X1 _7024_ (.A1(_2662_),
    .A2(_2664_),
    .ZN(_2665_));
 NAND2_X1 _7025_ (.A1(\aso.z0[1] ),
    .A2(_2306_),
    .ZN(_2666_));
 OAI21_X1 _7026_ (.A(_2662_),
    .B1(_2665_),
    .B2(_2666_),
    .ZN(_2667_));
 AOI21_X1 _7027_ (.A(_2587_),
    .B1(_2306_),
    .B2(\aso.z0[2] ),
    .ZN(_2668_));
 NOR2_X1 _7028_ (.A1(_2588_),
    .A2(_2668_),
    .ZN(_2669_));
 XNOR2_X1 _7029_ (.A(_2667_),
    .B(_2669_),
    .ZN(_2670_));
 NOR2_X1 _7030_ (.A1(_2661_),
    .A2(_2670_),
    .ZN(_2671_));
 AOI21_X1 _7031_ (.A(_2671_),
    .B1(_2669_),
    .B2(_2667_),
    .ZN(_2672_));
 XNOR2_X1 _7032_ (.A(_2595_),
    .B(_2596_),
    .ZN(_2673_));
 XNOR2_X1 _7033_ (.A(_2672_),
    .B(_2673_),
    .ZN(_2674_));
 NOR2_X1 _7034_ (.A1(_2659_),
    .A2(_2674_),
    .ZN(_2675_));
 NOR2_X1 _7035_ (.A1(_2672_),
    .A2(_2673_),
    .ZN(_2676_));
 OAI21_X1 _7036_ (.A(_2658_),
    .B1(_2675_),
    .B2(_2676_),
    .ZN(_2677_));
 OR3_X1 _7037_ (.A1(_2676_),
    .A2(_2675_),
    .A3(_2658_),
    .ZN(_2678_));
 AND2_X1 _7038_ (.A1(_2677_),
    .A2(_2678_),
    .ZN(_2679_));
 NAND2_X1 _7039_ (.A1(_2656_),
    .A2(_2679_),
    .ZN(_2680_));
 AOI21_X1 _7040_ (.A(_2636_),
    .B1(_2680_),
    .B2(_2677_),
    .ZN(_2681_));
 OR2_X1 _7041_ (.A1(_2639_),
    .A2(_2655_),
    .ZN(_2682_));
 OAI21_X1 _7042_ (.A(_2682_),
    .B1(_2654_),
    .B2(_2641_),
    .ZN(_2683_));
 NAND2_X1 _7043_ (.A1(_2677_),
    .A2(_2680_),
    .ZN(_2684_));
 XOR2_X1 _7044_ (.A(_2684_),
    .B(_2636_),
    .Z(_2685_));
 INV_X1 _7045_ (.A(_2685_),
    .ZN(_2686_));
 AOI21_X1 _7046_ (.A(_2681_),
    .B1(_2683_),
    .B2(_2686_),
    .ZN(_2687_));
 XNOR2_X1 _7047_ (.A(_2631_),
    .B(_2632_),
    .ZN(_2688_));
 NOR2_X1 _7048_ (.A1(_2687_),
    .A2(_2688_),
    .ZN(_2689_));
 XOR2_X1 _7049_ (.A(_2687_),
    .B(_2688_),
    .Z(_2690_));
 XOR2_X1 _7050_ (.A(_2659_),
    .B(_2674_),
    .Z(_2691_));
 INV_X1 _7051_ (.A(_2614_),
    .ZN(_2692_));
 OR3_X1 _7052_ (.A1(_0020_),
    .A2(_2692_),
    .A3(_2651_),
    .ZN(_2693_));
 OAI22_X1 _7053_ (.A1(_0020_),
    .A2(_2613_),
    .B1(_2692_),
    .B2(_2273_),
    .ZN(_2694_));
 AND2_X1 _7054_ (.A1(_2693_),
    .A2(_2694_),
    .ZN(_2695_));
 NAND3_X1 _7055_ (.A1(\aso.z0[8] ),
    .A2(_2637_),
    .A3(_2695_),
    .ZN(_2696_));
 NAND2_X1 _7056_ (.A1(_2693_),
    .A2(_2696_),
    .ZN(_2697_));
 INV_X1 _7057_ (.A(_2652_),
    .ZN(_2698_));
 OAI21_X1 _7058_ (.A(_2698_),
    .B1(_2650_),
    .B2(_2529_),
    .ZN(_2699_));
 XOR2_X1 _7059_ (.A(_2651_),
    .B(_2699_),
    .Z(_2700_));
 NAND2_X1 _7060_ (.A1(\aso.z0[4] ),
    .A2(_2449_),
    .ZN(_2701_));
 XOR2_X1 _7061_ (.A(_2480_),
    .B(_2701_),
    .Z(_2702_));
 NAND3_X1 _7062_ (.A1(\aso.z0[5] ),
    .A2(_2492_),
    .A3(_2702_),
    .ZN(_2703_));
 OAI21_X1 _7063_ (.A(_2703_),
    .B1(_2701_),
    .B2(_2480_),
    .ZN(_2704_));
 XOR2_X1 _7064_ (.A(_2700_),
    .B(_2704_),
    .Z(_2705_));
 XOR2_X1 _7065_ (.A(_2697_),
    .B(_2705_),
    .Z(_2706_));
 NAND4_X1 _7066_ (.A1(\aso.z0[2] ),
    .A2(_2501_),
    .A3(_2404_),
    .A4(_2449_),
    .ZN(_2707_));
 OAI22_X1 _7067_ (.A1(_2277_),
    .A2(_2437_),
    .B1(_2531_),
    .B2(_0011_),
    .ZN(_2708_));
 NAND2_X1 _7068_ (.A1(_2707_),
    .A2(_2708_),
    .ZN(_2709_));
 NAND2_X1 _7069_ (.A1(\aso.z0[1] ),
    .A2(_2342_),
    .ZN(_2710_));
 OAI21_X1 _7070_ (.A(_2707_),
    .B1(_2709_),
    .B2(_2710_),
    .ZN(_2711_));
 XOR2_X1 _7071_ (.A(_2665_),
    .B(_2666_),
    .Z(_2712_));
 XNOR2_X1 _7072_ (.A(_2711_),
    .B(_2712_),
    .ZN(_2713_));
 INV_X1 _7073_ (.A(_2713_),
    .ZN(_2714_));
 XNOR2_X1 _7074_ (.A(_2650_),
    .B(_2702_),
    .ZN(_2715_));
 AOI22_X1 _7075_ (.A1(_2711_),
    .A2(_2712_),
    .B1(_2714_),
    .B2(_2715_),
    .ZN(_2716_));
 XNOR2_X1 _7076_ (.A(_2661_),
    .B(_2670_),
    .ZN(_2717_));
 XOR2_X1 _7077_ (.A(_2716_),
    .B(_2717_),
    .Z(_2718_));
 AND2_X1 _7078_ (.A1(_2706_),
    .A2(_2718_),
    .ZN(_2719_));
 NOR2_X1 _7079_ (.A1(_2716_),
    .A2(_2717_),
    .ZN(_2720_));
 OAI21_X1 _7080_ (.A(_2691_),
    .B1(_2719_),
    .B2(_2720_),
    .ZN(_2721_));
 INV_X1 _7081_ (.A(_2721_),
    .ZN(_2722_));
 NAND2_X1 _7082_ (.A1(\aso.z0[8] ),
    .A2(_2637_),
    .ZN(_2723_));
 XOR2_X1 _7083_ (.A(\aso.z0[0] ),
    .B(\aso.z4[0] ),
    .Z(_2724_));
 OR2_X1 _7084_ (.A1(_0010_),
    .A2(_2724_),
    .ZN(_2725_));
 AOI22_X1 _7085_ (.A1(\aso.z0[8] ),
    .A2(_2614_),
    .B1(_2637_),
    .B2(\aso.z0[9] ),
    .ZN(_2726_));
 OAI22_X1 _7086_ (.A1(_2638_),
    .A2(_2723_),
    .B1(_2725_),
    .B2(_2726_),
    .ZN(_2727_));
 OAI21_X1 _7087_ (.A(_2638_),
    .B1(_2637_),
    .B2(_0010_),
    .ZN(_2728_));
 NAND2_X1 _7088_ (.A1(_2639_),
    .A2(_2728_),
    .ZN(_2729_));
 AND2_X1 _7089_ (.A1(_2700_),
    .A2(_2704_),
    .ZN(_2730_));
 AOI21_X1 _7090_ (.A(_2730_),
    .B1(_2705_),
    .B2(_2697_),
    .ZN(_2731_));
 XOR2_X1 _7091_ (.A(_2729_),
    .B(_2731_),
    .Z(_2732_));
 XOR2_X1 _7092_ (.A(_2727_),
    .B(_2732_),
    .Z(_2733_));
 NOR3_X1 _7093_ (.A1(_2720_),
    .A2(_2719_),
    .A3(_2691_),
    .ZN(_2734_));
 NOR2_X1 _7094_ (.A1(_2722_),
    .A2(_2734_),
    .ZN(_2735_));
 AOI21_X1 _7095_ (.A(_2722_),
    .B1(_2733_),
    .B2(_2735_),
    .ZN(_2736_));
 XNOR2_X1 _7096_ (.A(_2656_),
    .B(_2679_),
    .ZN(_2737_));
 NOR2_X1 _7097_ (.A1(_2736_),
    .A2(_2737_),
    .ZN(_2738_));
 NOR2_X1 _7098_ (.A1(_2729_),
    .A2(_2731_),
    .ZN(_2739_));
 AOI21_X1 _7099_ (.A(_2739_),
    .B1(_2732_),
    .B2(_2727_),
    .ZN(_2740_));
 INV_X1 _7100_ (.A(_2740_),
    .ZN(_2741_));
 XOR2_X1 _7101_ (.A(_2736_),
    .B(_2737_),
    .Z(_2742_));
 AOI21_X1 _7102_ (.A(_2738_),
    .B1(_2741_),
    .B2(_2742_),
    .ZN(_2743_));
 XOR2_X1 _7103_ (.A(_2683_),
    .B(_2685_),
    .Z(_2744_));
 XOR2_X1 _7104_ (.A(_2743_),
    .B(_2744_),
    .Z(_2745_));
 XOR2_X1 _7105_ (.A(_2733_),
    .B(_2735_),
    .Z(_2746_));
 NOR2_X1 _7106_ (.A1(_2638_),
    .A2(_2723_),
    .ZN(_2747_));
 NOR2_X1 _7107_ (.A1(_2747_),
    .A2(_2726_),
    .ZN(_2748_));
 XOR2_X1 _7108_ (.A(_2725_),
    .B(_2748_),
    .Z(_2749_));
 XOR2_X1 _7109_ (.A(_2695_),
    .B(_2723_),
    .Z(_2750_));
 NAND2_X1 _7110_ (.A1(\aso.z0[0] ),
    .A2(_2306_),
    .ZN(_2751_));
 NAND2_X1 _7111_ (.A1(\aso.z0[4] ),
    .A2(_2492_),
    .ZN(_2752_));
 XOR2_X1 _7112_ (.A(_2751_),
    .B(_2752_),
    .Z(_2753_));
 NAND3_X1 _7113_ (.A1(\aso.z0[5] ),
    .A2(_2566_),
    .A3(_2753_),
    .ZN(_2754_));
 OR2_X1 _7114_ (.A1(_2751_),
    .A2(_2752_),
    .ZN(_2755_));
 AOI21_X1 _7115_ (.A(_2750_),
    .B1(_2754_),
    .B2(_2755_),
    .ZN(_2756_));
 AND3_X1 _7116_ (.A1(_2755_),
    .A2(_2754_),
    .A3(_2750_),
    .ZN(_2757_));
 OR2_X1 _7117_ (.A1(_2756_),
    .A2(_2757_),
    .ZN(_2758_));
 INV_X1 _7118_ (.A(_2758_),
    .ZN(_2759_));
 INV_X1 _7119_ (.A(_2637_),
    .ZN(_2760_));
 OR4_X1 _7120_ (.A1(_2273_),
    .A2(_0020_),
    .A3(_2692_),
    .A4(_2760_),
    .ZN(_2761_));
 OAI22_X1 _7121_ (.A1(_0020_),
    .A2(_2692_),
    .B1(_2760_),
    .B2(_2273_),
    .ZN(_2762_));
 NAND2_X1 _7122_ (.A1(_2761_),
    .A2(_2762_),
    .ZN(_2763_));
 NAND2_X1 _7123_ (.A1(\aso.z0[8] ),
    .A2(_2724_),
    .ZN(_2764_));
 OAI21_X1 _7124_ (.A(_2761_),
    .B1(_2763_),
    .B2(_2764_),
    .ZN(_2765_));
 AOI21_X1 _7125_ (.A(_2756_),
    .B1(_2759_),
    .B2(_2765_),
    .ZN(_2766_));
 XOR2_X1 _7126_ (.A(_2749_),
    .B(_2766_),
    .Z(_2767_));
 NOR2_X1 _7127_ (.A1(_0011_),
    .A2(_2565_),
    .ZN(_2768_));
 NAND3_X1 _7128_ (.A1(\aso.z0[2] ),
    .A2(_2449_),
    .A3(_2768_),
    .ZN(_2769_));
 OAI22_X1 _7129_ (.A1(_2277_),
    .A2(_2531_),
    .B1(_2565_),
    .B2(_0011_),
    .ZN(_2770_));
 AND2_X1 _7130_ (.A1(_2769_),
    .A2(_2770_),
    .ZN(_2771_));
 AND3_X1 _7131_ (.A1(\aso.z0[1] ),
    .A2(_2404_),
    .A3(_2771_),
    .ZN(_2772_));
 INV_X1 _7132_ (.A(_2772_),
    .ZN(_2773_));
 NAND2_X1 _7133_ (.A1(_2769_),
    .A2(_2773_),
    .ZN(_2774_));
 XNOR2_X1 _7134_ (.A(_2709_),
    .B(_2710_),
    .ZN(_2775_));
 XNOR2_X1 _7135_ (.A(_2774_),
    .B(_2775_),
    .ZN(_2776_));
 NAND2_X1 _7136_ (.A1(\aso.z0[5] ),
    .A2(_2566_),
    .ZN(_2777_));
 XNOR2_X1 _7137_ (.A(_2777_),
    .B(_2753_),
    .ZN(_2778_));
 NAND2_X1 _7138_ (.A1(_2776_),
    .A2(_2778_),
    .ZN(_2779_));
 INV_X1 _7139_ (.A(_2774_),
    .ZN(_2780_));
 OAI21_X1 _7140_ (.A(_2779_),
    .B1(_2775_),
    .B2(_2780_),
    .ZN(_2781_));
 XNOR2_X1 _7141_ (.A(_2713_),
    .B(_2715_),
    .ZN(_2782_));
 NAND2_X1 _7142_ (.A1(_2781_),
    .A2(_2782_),
    .ZN(_2783_));
 XOR2_X1 _7143_ (.A(_2781_),
    .B(_2782_),
    .Z(_2784_));
 XNOR2_X1 _7144_ (.A(_2765_),
    .B(_2758_),
    .ZN(_2785_));
 NAND2_X1 _7145_ (.A1(_2784_),
    .A2(_2785_),
    .ZN(_2786_));
 NAND2_X1 _7146_ (.A1(_2783_),
    .A2(_2786_),
    .ZN(_2787_));
 XOR2_X1 _7147_ (.A(_2706_),
    .B(_2718_),
    .Z(_2788_));
 XOR2_X1 _7148_ (.A(_2787_),
    .B(_2788_),
    .Z(_2789_));
 AND2_X1 _7149_ (.A1(_2767_),
    .A2(_2789_),
    .ZN(_2790_));
 AND2_X1 _7150_ (.A1(_2787_),
    .A2(_2788_),
    .ZN(_2791_));
 OAI21_X1 _7151_ (.A(_2746_),
    .B1(_2790_),
    .B2(_2791_),
    .ZN(_2792_));
 NOR2_X1 _7152_ (.A1(_2749_),
    .A2(_2766_),
    .ZN(_2793_));
 OR3_X1 _7153_ (.A1(_2791_),
    .A2(_2790_),
    .A3(_2746_),
    .ZN(_2794_));
 AND2_X1 _7154_ (.A1(_2792_),
    .A2(_2794_),
    .ZN(_2795_));
 NAND2_X1 _7155_ (.A1(_2793_),
    .A2(_2795_),
    .ZN(_2796_));
 NAND2_X1 _7156_ (.A1(_2792_),
    .A2(_2796_),
    .ZN(_2797_));
 XNOR2_X1 _7157_ (.A(_2740_),
    .B(_2742_),
    .ZN(_2798_));
 NAND2_X1 _7158_ (.A1(_2797_),
    .A2(_2798_),
    .ZN(_2799_));
 XOR2_X1 _7159_ (.A(_2797_),
    .B(_2798_),
    .Z(_2800_));
 XOR2_X1 _7160_ (.A(_2767_),
    .B(_2789_),
    .Z(_2801_));
 XNOR2_X1 _7161_ (.A(_2784_),
    .B(_2785_),
    .ZN(_2802_));
 XOR2_X1 _7162_ (.A(_2776_),
    .B(_2778_),
    .Z(_2803_));
 NAND3_X1 _7163_ (.A1(\aso.z0[2] ),
    .A2(_2566_),
    .A3(_2768_),
    .ZN(_2804_));
 OAI22_X1 _7164_ (.A1(_2277_),
    .A2(_2565_),
    .B1(_2613_),
    .B2(_0011_),
    .ZN(_2805_));
 NAND4_X1 _7165_ (.A1(\aso.z0[1] ),
    .A2(_2449_),
    .A3(_2804_),
    .A4(_2805_),
    .ZN(_2806_));
 NAND2_X1 _7166_ (.A1(_2804_),
    .A2(_2806_),
    .ZN(_2807_));
 AOI21_X1 _7167_ (.A(_2771_),
    .B1(_2404_),
    .B2(\aso.z0[1] ),
    .ZN(_2808_));
 NOR2_X1 _7168_ (.A1(_2772_),
    .A2(_2808_),
    .ZN(_2809_));
 XNOR2_X1 _7169_ (.A(_2807_),
    .B(_2809_),
    .ZN(_2810_));
 NAND2_X1 _7170_ (.A1(\aso.z0[5] ),
    .A2(_2614_),
    .ZN(_2811_));
 NAND2_X1 _7171_ (.A1(\aso.z0[4] ),
    .A2(_2566_),
    .ZN(_2812_));
 XOR2_X1 _7172_ (.A(_2605_),
    .B(_2812_),
    .Z(_2813_));
 XNOR2_X1 _7173_ (.A(_2811_),
    .B(_2813_),
    .ZN(_2814_));
 INV_X1 _7174_ (.A(_2814_),
    .ZN(_2815_));
 NOR2_X1 _7175_ (.A1(_2810_),
    .A2(_2815_),
    .ZN(_2816_));
 AND2_X1 _7176_ (.A1(_2807_),
    .A2(_2809_),
    .ZN(_2817_));
 OAI21_X1 _7177_ (.A(_2803_),
    .B1(_2816_),
    .B2(_2817_),
    .ZN(_2818_));
 OR3_X1 _7178_ (.A1(_2817_),
    .A2(_2816_),
    .A3(_2803_),
    .ZN(_2819_));
 AND2_X1 _7179_ (.A1(_2818_),
    .A2(_2819_),
    .ZN(_2820_));
 NAND2_X1 _7180_ (.A1(\aso.z0[7] ),
    .A2(_2724_),
    .ZN(_2821_));
 NAND2_X1 _7181_ (.A1(\aso.z0[6] ),
    .A2(_2637_),
    .ZN(_2822_));
 NOR2_X1 _7182_ (.A1(_2821_),
    .A2(_2822_),
    .ZN(_2823_));
 XOR2_X1 _7183_ (.A(_2763_),
    .B(_2764_),
    .Z(_2824_));
 NAND3_X1 _7184_ (.A1(\aso.z0[5] ),
    .A2(_2614_),
    .A3(_2813_),
    .ZN(_2825_));
 OAI21_X1 _7185_ (.A(_2825_),
    .B1(_2812_),
    .B2(_2605_),
    .ZN(_2826_));
 XOR2_X1 _7186_ (.A(_2824_),
    .B(_2826_),
    .Z(_2827_));
 XOR2_X1 _7187_ (.A(_2823_),
    .B(_2827_),
    .Z(_2828_));
 NAND2_X1 _7188_ (.A1(_2820_),
    .A2(_2828_),
    .ZN(_2829_));
 AOI21_X1 _7189_ (.A(_2802_),
    .B1(_2829_),
    .B2(_2818_),
    .ZN(_2830_));
 AND3_X1 _7190_ (.A1(_2818_),
    .A2(_2829_),
    .A3(_2802_),
    .ZN(_2831_));
 NOR2_X1 _7191_ (.A1(_2830_),
    .A2(_2831_),
    .ZN(_2832_));
 NAND2_X1 _7192_ (.A1(\aso.z0[9] ),
    .A2(_2724_),
    .ZN(_2833_));
 AOI22_X1 _7193_ (.A1(_2824_),
    .A2(_2826_),
    .B1(_2827_),
    .B2(_2823_),
    .ZN(_2834_));
 XOR2_X1 _7194_ (.A(_2833_),
    .B(_2834_),
    .Z(_2835_));
 AND2_X1 _7195_ (.A1(_2832_),
    .A2(_2835_),
    .ZN(_2836_));
 OAI21_X1 _7196_ (.A(_2801_),
    .B1(_2836_),
    .B2(_2830_),
    .ZN(_2837_));
 INV_X1 _7197_ (.A(_2837_),
    .ZN(_2838_));
 NOR3_X1 _7198_ (.A1(_2830_),
    .A2(_2836_),
    .A3(_2801_),
    .ZN(_2839_));
 NOR2_X1 _7199_ (.A1(_2838_),
    .A2(_2839_),
    .ZN(_2840_));
 NOR2_X1 _7200_ (.A1(_2833_),
    .A2(_2834_),
    .ZN(_2841_));
 AOI21_X1 _7201_ (.A(_2838_),
    .B1(_2840_),
    .B2(_2841_),
    .ZN(_2842_));
 XNOR2_X1 _7202_ (.A(_2793_),
    .B(_2795_),
    .ZN(_2843_));
 NOR2_X1 _7203_ (.A1(_2842_),
    .A2(_2843_),
    .ZN(_2844_));
 XNOR2_X1 _7204_ (.A(_2842_),
    .B(_2843_),
    .ZN(_2845_));
 XNOR2_X1 _7205_ (.A(_2820_),
    .B(_2828_),
    .ZN(_2846_));
 XNOR2_X1 _7206_ (.A(_2810_),
    .B(_2814_),
    .ZN(_2847_));
 NOR2_X1 _7207_ (.A1(_0011_),
    .A2(_2692_),
    .ZN(_2848_));
 NAND3_X1 _7208_ (.A1(\aso.z0[2] ),
    .A2(_2566_),
    .A3(_2848_),
    .ZN(_2849_));
 OAI22_X1 _7209_ (.A1(_2277_),
    .A2(_2613_),
    .B1(_2692_),
    .B2(_0011_),
    .ZN(_2850_));
 AND2_X1 _7210_ (.A1(_2849_),
    .A2(_2850_),
    .ZN(_2851_));
 NAND3_X1 _7211_ (.A1(\aso.z0[1] ),
    .A2(_2492_),
    .A3(_2851_),
    .ZN(_2852_));
 NAND2_X1 _7212_ (.A1(_2849_),
    .A2(_2852_),
    .ZN(_2853_));
 NAND2_X1 _7213_ (.A1(_2804_),
    .A2(_2805_),
    .ZN(_2854_));
 OAI21_X1 _7214_ (.A(_2854_),
    .B1(_2531_),
    .B2(_2278_),
    .ZN(_2855_));
 NAND2_X1 _7215_ (.A1(_2806_),
    .A2(_2855_),
    .ZN(_2856_));
 XNOR2_X1 _7216_ (.A(_2853_),
    .B(_2856_),
    .ZN(_2857_));
 NAND2_X1 _7217_ (.A1(\aso.z0[5] ),
    .A2(_2637_),
    .ZN(_2858_));
 NAND4_X1 _7218_ (.A1(\aso.z0[4] ),
    .A2(\aso.z0[0] ),
    .A3(_2404_),
    .A4(_2614_),
    .ZN(_2859_));
 OAI22_X1 _7219_ (.A1(_2280_),
    .A2(_2437_),
    .B1(_2692_),
    .B2(_2275_),
    .ZN(_2860_));
 AND2_X1 _7220_ (.A1(_2859_),
    .A2(_2860_),
    .ZN(_2861_));
 XNOR2_X1 _7221_ (.A(_2858_),
    .B(_2861_),
    .ZN(_2862_));
 AND2_X1 _7222_ (.A1(_2857_),
    .A2(_2862_),
    .ZN(_2863_));
 AOI21_X1 _7223_ (.A(_2856_),
    .B1(_2852_),
    .B2(_2849_),
    .ZN(_2864_));
 OAI21_X1 _7224_ (.A(_2847_),
    .B1(_2863_),
    .B2(_2864_),
    .ZN(_2865_));
 OR3_X1 _7225_ (.A1(_2864_),
    .A2(_2863_),
    .A3(_2847_),
    .ZN(_2866_));
 AND2_X1 _7226_ (.A1(_2865_),
    .A2(_2866_),
    .ZN(_2867_));
 XNOR2_X1 _7227_ (.A(_2821_),
    .B(_2822_),
    .ZN(_2868_));
 NAND3_X1 _7228_ (.A1(\aso.z0[5] ),
    .A2(_2637_),
    .A3(_2861_),
    .ZN(_2869_));
 AOI21_X1 _7229_ (.A(_2868_),
    .B1(_2869_),
    .B2(_2859_),
    .ZN(_2870_));
 AND3_X1 _7230_ (.A1(_2859_),
    .A2(_2869_),
    .A3(_2868_),
    .ZN(_2871_));
 NOR2_X1 _7231_ (.A1(_2870_),
    .A2(_2871_),
    .ZN(_2872_));
 NAND2_X1 _7232_ (.A1(_2867_),
    .A2(_2872_),
    .ZN(_2873_));
 AOI21_X1 _7233_ (.A(_2846_),
    .B1(_2873_),
    .B2(_2865_),
    .ZN(_2874_));
 AND3_X1 _7234_ (.A1(_2865_),
    .A2(_2873_),
    .A3(_2846_),
    .ZN(_2875_));
 NOR2_X1 _7235_ (.A1(_2874_),
    .A2(_2875_),
    .ZN(_2876_));
 AOI21_X1 _7236_ (.A(_2874_),
    .B1(_2876_),
    .B2(_2870_),
    .ZN(_2877_));
 XNOR2_X1 _7237_ (.A(_2832_),
    .B(_2835_),
    .ZN(_2878_));
 XNOR2_X1 _7238_ (.A(_2841_),
    .B(_2840_),
    .ZN(_2879_));
 OR3_X1 _7239_ (.A1(_2877_),
    .A2(_2878_),
    .A3(_2879_),
    .ZN(_2880_));
 NOR2_X1 _7240_ (.A1(_2877_),
    .A2(_2878_),
    .ZN(_2881_));
 XNOR2_X1 _7241_ (.A(_2881_),
    .B(_2879_),
    .ZN(_2882_));
 NAND4_X1 _7242_ (.A1(\aso.z0[4] ),
    .A2(\aso.z0[0] ),
    .A3(_2449_),
    .A4(_2637_),
    .ZN(_2883_));
 OAI22_X1 _7243_ (.A1(_2280_),
    .A2(_2531_),
    .B1(_2760_),
    .B2(_2275_),
    .ZN(_2884_));
 AND2_X1 _7244_ (.A1(_2883_),
    .A2(_2884_),
    .ZN(_2885_));
 NAND3_X1 _7245_ (.A1(\aso.z0[5] ),
    .A2(_2724_),
    .A3(_2885_),
    .ZN(_2886_));
 NAND2_X1 _7246_ (.A1(_2883_),
    .A2(_2886_),
    .ZN(_2887_));
 AND3_X1 _7247_ (.A1(\aso.z0[6] ),
    .A2(_2724_),
    .A3(_2887_),
    .ZN(_2888_));
 XOR2_X1 _7248_ (.A(_2857_),
    .B(_2862_),
    .Z(_2889_));
 NOR2_X1 _7249_ (.A1(_2277_),
    .A2(_2760_),
    .ZN(_2890_));
 NAND2_X1 _7250_ (.A1(_2848_),
    .A2(_2890_),
    .ZN(_2891_));
 AOI22_X1 _7251_ (.A1(\aso.z0[2] ),
    .A2(_2614_),
    .B1(_2637_),
    .B2(_2501_),
    .ZN(_2892_));
 AOI21_X1 _7252_ (.A(_2892_),
    .B1(_2890_),
    .B2(_2848_),
    .ZN(_2893_));
 NAND3_X1 _7253_ (.A1(\aso.z0[1] ),
    .A2(_2566_),
    .A3(_2893_),
    .ZN(_2894_));
 NAND2_X1 _7254_ (.A1(_2891_),
    .A2(_2894_),
    .ZN(_2895_));
 NAND2_X1 _7255_ (.A1(\aso.z0[1] ),
    .A2(_2492_),
    .ZN(_2896_));
 XOR2_X1 _7256_ (.A(_2851_),
    .B(_2896_),
    .Z(_2897_));
 XNOR2_X1 _7257_ (.A(_2895_),
    .B(_2897_),
    .ZN(_2898_));
 NAND2_X1 _7258_ (.A1(\aso.z0[5] ),
    .A2(_2724_),
    .ZN(_2899_));
 XNOR2_X1 _7259_ (.A(_2899_),
    .B(_2885_),
    .ZN(_2900_));
 AND2_X1 _7260_ (.A1(_2898_),
    .A2(_2900_),
    .ZN(_2901_));
 AOI21_X1 _7261_ (.A(_2897_),
    .B1(_2894_),
    .B2(_2891_),
    .ZN(_2902_));
 OAI21_X1 _7262_ (.A(_2889_),
    .B1(_2901_),
    .B2(_2902_),
    .ZN(_2903_));
 INV_X1 _7263_ (.A(_2903_),
    .ZN(_2904_));
 NOR3_X1 _7264_ (.A1(_2902_),
    .A2(_2901_),
    .A3(_2889_),
    .ZN(_2905_));
 NOR2_X1 _7265_ (.A1(_2904_),
    .A2(_2905_),
    .ZN(_2906_));
 AOI21_X1 _7266_ (.A(_2887_),
    .B1(_2724_),
    .B2(\aso.z0[6] ),
    .ZN(_2907_));
 NOR2_X1 _7267_ (.A1(_2907_),
    .A2(_2888_),
    .ZN(_2908_));
 AOI21_X1 _7268_ (.A(_2904_),
    .B1(_2906_),
    .B2(_2908_),
    .ZN(_2909_));
 XNOR2_X1 _7269_ (.A(_2867_),
    .B(_2872_),
    .ZN(_2910_));
 XOR2_X1 _7270_ (.A(_2909_),
    .B(_2910_),
    .Z(_2911_));
 NAND2_X1 _7271_ (.A1(_2888_),
    .A2(_2911_),
    .ZN(_2912_));
 OAI21_X1 _7272_ (.A(_2912_),
    .B1(_2910_),
    .B2(_2909_),
    .ZN(_2913_));
 XOR2_X1 _7273_ (.A(_2870_),
    .B(_2876_),
    .Z(_2914_));
 AND2_X1 _7274_ (.A1(_2913_),
    .A2(_2914_),
    .ZN(_2915_));
 XOR2_X1 _7275_ (.A(_2877_),
    .B(_2878_),
    .Z(_2916_));
 NAND2_X1 _7276_ (.A1(_2915_),
    .A2(_2916_),
    .ZN(_2917_));
 XNOR2_X1 _7277_ (.A(_2915_),
    .B(_2916_),
    .ZN(_2918_));
 XOR2_X1 _7278_ (.A(_2888_),
    .B(_2911_),
    .Z(_2919_));
 INV_X1 _7279_ (.A(_2724_),
    .ZN(_2920_));
 NOR2_X1 _7280_ (.A1(_0011_),
    .A2(_2920_),
    .ZN(_2921_));
 XOR2_X1 _7281_ (.A(_2890_),
    .B(_2921_),
    .Z(_2922_));
 AND3_X1 _7282_ (.A1(\aso.z0[1] ),
    .A2(_2614_),
    .A3(_2922_),
    .ZN(_2923_));
 AOI21_X1 _7283_ (.A(_2923_),
    .B1(_2921_),
    .B2(_2890_),
    .ZN(_2924_));
 NAND2_X1 _7284_ (.A1(\aso.z0[1] ),
    .A2(_2566_),
    .ZN(_2925_));
 XOR2_X1 _7285_ (.A(_2893_),
    .B(_2925_),
    .Z(_2926_));
 XNOR2_X1 _7286_ (.A(_2924_),
    .B(_2926_),
    .ZN(_2927_));
 NOR3_X1 _7287_ (.A1(_2280_),
    .A2(\aso.z4[0] ),
    .A3(_2752_),
    .ZN(_2928_));
 AOI22_X1 _7288_ (.A1(\aso.z0[0] ),
    .A2(_2492_),
    .B1(_2724_),
    .B2(\aso.z0[4] ),
    .ZN(_2929_));
 NOR2_X1 _7289_ (.A1(_2928_),
    .A2(_2929_),
    .ZN(_2930_));
 INV_X1 _7290_ (.A(_2930_),
    .ZN(_2931_));
 OAI22_X1 _7291_ (.A1(_2924_),
    .A2(_2926_),
    .B1(_2927_),
    .B2(_2931_),
    .ZN(_2932_));
 XOR2_X1 _7292_ (.A(_2898_),
    .B(_2900_),
    .Z(_2933_));
 XOR2_X1 _7293_ (.A(_2932_),
    .B(_2933_),
    .Z(_2934_));
 AOI22_X1 _7294_ (.A1(_2932_),
    .A2(_2933_),
    .B1(_2934_),
    .B2(_2928_),
    .ZN(_2935_));
 XNOR2_X1 _7295_ (.A(_2906_),
    .B(_2908_),
    .ZN(_2936_));
 NOR2_X1 _7296_ (.A1(_2935_),
    .A2(_2936_),
    .ZN(_2937_));
 AND2_X1 _7297_ (.A1(_2935_),
    .A2(_2936_),
    .ZN(_2938_));
 NOR2_X1 _7298_ (.A1(_2280_),
    .A2(_2613_),
    .ZN(_2939_));
 NAND4_X1 _7299_ (.A1(\aso.z0[2] ),
    .A2(\aso.z0[1] ),
    .A3(_2637_),
    .A4(_2724_),
    .ZN(_2940_));
 AOI21_X1 _7300_ (.A(_2922_),
    .B1(_2614_),
    .B2(\aso.z0[1] ),
    .ZN(_2941_));
 NOR2_X1 _7301_ (.A1(_2923_),
    .A2(_2941_),
    .ZN(_2942_));
 XNOR2_X1 _7302_ (.A(_2940_),
    .B(_2942_),
    .ZN(_2943_));
 XOR2_X1 _7303_ (.A(_2939_),
    .B(_2943_),
    .Z(_2944_));
 XOR2_X1 _7304_ (.A(_2927_),
    .B(_2930_),
    .Z(_2945_));
 NOR3_X1 _7305_ (.A1(_2923_),
    .A2(_2940_),
    .A3(_2941_),
    .ZN(_2946_));
 AOI21_X1 _7306_ (.A(_2946_),
    .B1(_2943_),
    .B2(_2939_),
    .ZN(_2947_));
 OAI21_X1 _7307_ (.A(_2944_),
    .B1(_2945_),
    .B2(_2947_),
    .ZN(_2948_));
 AOI21_X1 _7308_ (.A(_2948_),
    .B1(_2945_),
    .B2(_2947_),
    .ZN(_2949_));
 XOR2_X1 _7309_ (.A(_2928_),
    .B(_2934_),
    .Z(_2950_));
 OAI22_X1 _7310_ (.A1(_2278_),
    .A2(_2760_),
    .B1(_2920_),
    .B2(_2277_),
    .ZN(_2951_));
 AND2_X1 _7311_ (.A1(_2940_),
    .A2(_2951_),
    .ZN(_2952_));
 NAND3_X1 _7312_ (.A1(\aso.z0[0] ),
    .A2(_2614_),
    .A3(_2952_),
    .ZN(_2953_));
 INV_X1 _7313_ (.A(_2953_),
    .ZN(_2954_));
 AND2_X1 _7314_ (.A1(_2950_),
    .A2(_2954_),
    .ZN(_2955_));
 NOR2_X1 _7315_ (.A1(_2614_),
    .A2(_2952_),
    .ZN(_2956_));
 NAND4_X1 _7316_ (.A1(\aso.z0[1] ),
    .A2(\aso.z0[0] ),
    .A3(_2637_),
    .A4(_2724_),
    .ZN(_2957_));
 NOR3_X1 _7317_ (.A1(_2954_),
    .A2(_2956_),
    .A3(_2957_),
    .ZN(_2958_));
 NOR2_X1 _7318_ (.A1(_2947_),
    .A2(_2945_),
    .ZN(_2959_));
 XOR2_X1 _7319_ (.A(_2950_),
    .B(_2959_),
    .Z(_2960_));
 AND2_X1 _7320_ (.A1(_2944_),
    .A2(_2954_),
    .ZN(_2961_));
 OAI221_X1 _7321_ (.A(_2949_),
    .B1(_2955_),
    .B2(_2958_),
    .C1(_2960_),
    .C2(_2961_),
    .ZN(_2963_));
 NAND2_X1 _7322_ (.A1(_2950_),
    .A2(_2959_),
    .ZN(_2964_));
 AOI211_X1 _7323_ (.A(_2937_),
    .B(_2938_),
    .C1(_2963_),
    .C2(_2964_),
    .ZN(_2965_));
 OAI21_X1 _7324_ (.A(_2919_),
    .B1(_2965_),
    .B2(_2937_),
    .ZN(_2966_));
 NOR2_X1 _7325_ (.A1(_2915_),
    .A2(_2966_),
    .ZN(_2967_));
 OAI21_X1 _7326_ (.A(_2967_),
    .B1(_2914_),
    .B2(_2913_),
    .ZN(_2968_));
 OAI21_X1 _7327_ (.A(_2917_),
    .B1(_2918_),
    .B2(_2968_),
    .ZN(_2969_));
 NAND2_X1 _7328_ (.A1(_2882_),
    .A2(_2969_),
    .ZN(_2970_));
 AOI21_X1 _7329_ (.A(_2845_),
    .B1(_2880_),
    .B2(_2970_),
    .ZN(_2971_));
 OAI21_X1 _7330_ (.A(_2800_),
    .B1(_2844_),
    .B2(_2971_),
    .ZN(_2972_));
 NAND2_X1 _7331_ (.A1(_2799_),
    .A2(_2972_),
    .ZN(_2974_));
 NAND2_X1 _7332_ (.A1(_2745_),
    .A2(_2974_),
    .ZN(_2975_));
 OAI21_X1 _7333_ (.A(_2975_),
    .B1(_2744_),
    .B2(_2743_),
    .ZN(_2976_));
 AOI21_X1 _7334_ (.A(_2689_),
    .B1(_2690_),
    .B2(_2976_),
    .ZN(_2977_));
 NOR2_X1 _7335_ (.A1(_2635_),
    .A2(_2977_),
    .ZN(_2978_));
 INV_X1 _7336_ (.A(_2634_),
    .ZN(_2979_));
 AOI21_X1 _7337_ (.A(_2978_),
    .B1(_2979_),
    .B2(_2633_),
    .ZN(_2980_));
 XOR2_X1 _7338_ (.A(_2581_),
    .B(_2583_),
    .Z(_2981_));
 NOR2_X1 _7339_ (.A1(_2980_),
    .A2(_2981_),
    .ZN(_2982_));
 AOI211_X1 _7340_ (.A(_2525_),
    .B(_2585_),
    .C1(_2982_),
    .C2(_2527_),
    .ZN(_2983_));
 XOR2_X1 _7341_ (.A(_2466_),
    .B(_2467_),
    .Z(_2985_));
 OR2_X1 _7342_ (.A1(_2983_),
    .A2(_2985_),
    .ZN(_2986_));
 NAND2_X1 _7343_ (.A1(_2469_),
    .A2(_2986_),
    .ZN(_2987_));
 XNOR2_X1 _7344_ (.A(_2424_),
    .B(_2987_),
    .ZN(_2988_));
 XNOR2_X1 _7345_ (.A(_2983_),
    .B(_2985_),
    .ZN(_2989_));
 NOR2_X1 _7346_ (.A1(_2584_),
    .A2(_2982_),
    .ZN(_2990_));
 XOR2_X1 _7347_ (.A(_2527_),
    .B(_2990_),
    .Z(_2991_));
 XOR2_X1 _7348_ (.A(_2980_),
    .B(_2981_),
    .Z(_2992_));
 XOR2_X1 _7349_ (.A(_2635_),
    .B(_2977_),
    .Z(_2993_));
 XOR2_X1 _7350_ (.A(_2690_),
    .B(_2976_),
    .Z(_2994_));
 NOR2_X1 _7351_ (.A1(_2844_),
    .A2(_2971_),
    .ZN(_2996_));
 XNOR2_X1 _7352_ (.A(_2800_),
    .B(_2996_),
    .ZN(_2997_));
 XNOR2_X1 _7353_ (.A(_2918_),
    .B(_2968_),
    .ZN(_2998_));
 XNOR2_X1 _7354_ (.A(_2882_),
    .B(_2969_),
    .ZN(_2999_));
 NOR2_X1 _7355_ (.A1(_2998_),
    .A2(_2999_),
    .ZN(_3000_));
 AND3_X1 _7356_ (.A1(_2845_),
    .A2(_2880_),
    .A3(_2970_),
    .ZN(_3001_));
 NOR2_X1 _7357_ (.A1(_2971_),
    .A2(_3001_),
    .ZN(_3002_));
 AND2_X1 _7358_ (.A1(_3000_),
    .A2(_3002_),
    .ZN(_3003_));
 AND2_X1 _7359_ (.A1(_2997_),
    .A2(_3003_),
    .ZN(_3004_));
 XOR2_X1 _7360_ (.A(_2745_),
    .B(_2974_),
    .Z(_3005_));
 AND2_X1 _7361_ (.A1(_3004_),
    .A2(_3005_),
    .ZN(_3007_));
 AND2_X1 _7362_ (.A1(_2994_),
    .A2(_3007_),
    .ZN(_3008_));
 AND2_X1 _7363_ (.A1(_2993_),
    .A2(_3008_),
    .ZN(_3009_));
 NAND2_X1 _7364_ (.A1(_2992_),
    .A2(_3009_),
    .ZN(_3010_));
 OR2_X1 _7365_ (.A1(_2991_),
    .A2(_3010_),
    .ZN(_3011_));
 NOR2_X1 _7366_ (.A1(_2989_),
    .A2(_3011_),
    .ZN(_3012_));
 OAI21_X1 _7367_ (.A(_2962_),
    .B1(_2988_),
    .B2(_3012_),
    .ZN(_3013_));
 AOI21_X1 _7368_ (.A(_3013_),
    .B1(_3012_),
    .B2(_2988_),
    .ZN(_0051_));
 AND2_X1 _7369_ (.A1(_2989_),
    .A2(_3011_),
    .ZN(_3014_));
 NOR3_X1 _7370_ (.A1(rst),
    .A2(_3012_),
    .A3(_3014_),
    .ZN(_0050_));
 NAND2_X1 _7371_ (.A1(_2962_),
    .A2(_3011_),
    .ZN(_3016_));
 AOI21_X1 _7372_ (.A(_3016_),
    .B1(_3010_),
    .B2(_2991_),
    .ZN(_0049_));
 OAI21_X1 _7373_ (.A(_2962_),
    .B1(_2992_),
    .B2(_3009_),
    .ZN(_3017_));
 AOI21_X1 _7374_ (.A(_3017_),
    .B1(_3009_),
    .B2(_2992_),
    .ZN(_0048_));
 NOR2_X1 _7375_ (.A1(_2993_),
    .A2(_3008_),
    .ZN(_3018_));
 NOR3_X1 _7376_ (.A1(rst),
    .A2(_3009_),
    .A3(_3018_),
    .ZN(_0047_));
 NOR2_X1 _7377_ (.A1(_2994_),
    .A2(_3007_),
    .ZN(_3019_));
 NOR3_X1 _7378_ (.A1(rst),
    .A2(_3008_),
    .A3(_3019_),
    .ZN(_0046_));
 NOR2_X1 _7379_ (.A1(_3004_),
    .A2(_3005_),
    .ZN(_3020_));
 NOR3_X1 _7380_ (.A1(rst),
    .A2(_3007_),
    .A3(_3020_),
    .ZN(_0045_));
 NOR2_X1 _7381_ (.A1(_2997_),
    .A2(_3003_),
    .ZN(_3022_));
 NOR3_X1 _7382_ (.A1(rst),
    .A2(_3004_),
    .A3(_3022_),
    .ZN(_0044_));
 NOR2_X1 _7383_ (.A1(_3000_),
    .A2(_3002_),
    .ZN(_3023_));
 NOR3_X1 _7384_ (.A1(rst),
    .A2(_3003_),
    .A3(_3023_),
    .ZN(_0043_));
 INV_X1 _7385_ (.A(_2469_),
    .ZN(_3024_));
 AOI21_X1 _7386_ (.A(_2421_),
    .B1(_2423_),
    .B2(_3024_),
    .ZN(_3025_));
 OAI21_X1 _7387_ (.A(_3025_),
    .B1(_2986_),
    .B2(_2424_),
    .ZN(_3026_));
 INV_X1 _7388_ (.A(_2388_),
    .ZN(_3027_));
 NOR2_X1 _7389_ (.A1(_2345_),
    .A2(_3027_),
    .ZN(_3028_));
 INV_X1 _7390_ (.A(_2387_),
    .ZN(_3029_));
 AOI21_X1 _7391_ (.A(_3028_),
    .B1(_3029_),
    .B2(_2369_),
    .ZN(_3031_));
 NOR2_X1 _7392_ (.A1(_2373_),
    .A2(_2375_),
    .ZN(_3032_));
 NOR2_X1 _7393_ (.A1(_2370_),
    .A2(_2376_),
    .ZN(_3033_));
 NOR2_X1 _7394_ (.A1(_3032_),
    .A2(_3033_),
    .ZN(_3034_));
 AOI21_X1 _7395_ (.A(_2384_),
    .B1(_2386_),
    .B2(_2377_),
    .ZN(_3035_));
 OR2_X1 _7396_ (.A1(_2350_),
    .A2(_2381_),
    .ZN(_3036_));
 NAND3_X1 _7397_ (.A1(_2350_),
    .A2(_2354_),
    .A3(_2381_),
    .ZN(_3037_));
 NAND2_X1 _7398_ (.A1(_3036_),
    .A2(_3037_),
    .ZN(_3038_));
 NAND3_X1 _7399_ (.A1(\aso.z0[9] ),
    .A2(_2318_),
    .A3(_2371_),
    .ZN(_3039_));
 OAI21_X1 _7400_ (.A(_2372_),
    .B1(_2318_),
    .B2(_2279_),
    .ZN(_3040_));
 INV_X1 _7401_ (.A(_3040_),
    .ZN(_3042_));
 NOR2_X1 _7402_ (.A1(_2374_),
    .A2(_2379_),
    .ZN(_3043_));
 XNOR2_X1 _7403_ (.A(_3042_),
    .B(_3043_),
    .ZN(_3044_));
 XNOR2_X1 _7404_ (.A(_3039_),
    .B(_3044_),
    .ZN(_3045_));
 XNOR2_X1 _7405_ (.A(_3038_),
    .B(_3045_),
    .ZN(_3046_));
 XNOR2_X1 _7406_ (.A(_3035_),
    .B(_3046_),
    .ZN(_3047_));
 XNOR2_X1 _7407_ (.A(_3034_),
    .B(_3047_),
    .ZN(_3048_));
 XOR2_X1 _7408_ (.A(_3031_),
    .B(_3048_),
    .Z(_3049_));
 NAND2_X1 _7409_ (.A1(_3026_),
    .A2(_3049_),
    .ZN(_3050_));
 OAI21_X1 _7410_ (.A(_3050_),
    .B1(_3048_),
    .B2(_3031_),
    .ZN(_3051_));
 NOR2_X1 _7411_ (.A1(_3035_),
    .A2(_3046_),
    .ZN(_3053_));
 NOR2_X1 _7412_ (.A1(_3034_),
    .A2(_3047_),
    .ZN(_3054_));
 NOR2_X1 _7413_ (.A1(_3053_),
    .A2(_3054_),
    .ZN(_3055_));
 OAI22_X1 _7414_ (.A1(_3042_),
    .A2(_3043_),
    .B1(_3044_),
    .B2(_3039_),
    .ZN(_3056_));
 OAI22_X1 _7415_ (.A1(_3039_),
    .A2(_3038_),
    .B1(_3044_),
    .B2(_3036_),
    .ZN(_3057_));
 INV_X1 _7416_ (.A(_3037_),
    .ZN(_3058_));
 AOI21_X1 _7417_ (.A(_3057_),
    .B1(_3044_),
    .B2(_3058_),
    .ZN(_3059_));
 XNOR2_X1 _7418_ (.A(_3056_),
    .B(_3059_),
    .ZN(_3060_));
 XNOR2_X1 _7419_ (.A(_3055_),
    .B(_3060_),
    .ZN(_3061_));
 NAND2_X1 _7420_ (.A1(_2988_),
    .A2(_3012_),
    .ZN(_3062_));
 XNOR2_X1 _7421_ (.A(_3026_),
    .B(_3049_),
    .ZN(_3064_));
 NOR2_X1 _7422_ (.A1(_3062_),
    .A2(_3064_),
    .ZN(_3065_));
 NOR2_X1 _7423_ (.A1(rst),
    .A2(_3065_),
    .ZN(_3066_));
 INV_X1 _7424_ (.A(_3066_),
    .ZN(_3067_));
 NOR3_X1 _7425_ (.A1(_3051_),
    .A2(_3061_),
    .A3(_3067_),
    .ZN(_0042_));
 AOI21_X1 _7426_ (.A(_3067_),
    .B1(_3064_),
    .B2(_3062_),
    .ZN(_0041_));
 AND2_X1 _7427_ (.A1(_2998_),
    .A2(_2999_),
    .ZN(_3068_));
 NOR3_X1 _7428_ (.A1(rst),
    .A2(_3000_),
    .A3(_3068_),
    .ZN(_0040_));
 DFF_X1 \aso.p[0]$_SDFF_PP0_  (.D(_0040_),
    .CK(clknet_4_4_0_clk),
    .Q(\aso.p[0] ),
    .QN(_3801_));
 DFF_X1 \aso.p[10]$_SDFF_PP0_  (.D(_0041_),
    .CK(clknet_4_14_0_clk),
    .Q(\aso.p[10] ),
    .QN(_3800_));
 DFF_X1 \aso.p[11]$_SDFF_PP0_  (.D(_0042_),
    .CK(clknet_4_15_0_clk),
    .Q(\aso.p[11] ),
    .QN(_3799_));
 DFF_X1 \aso.p[1]$_SDFF_PP0_  (.D(_0043_),
    .CK(clknet_4_10_0_clk),
    .Q(\aso.p[1] ),
    .QN(_3798_));
 DFF_X1 \aso.p[2]$_SDFF_PP0_  (.D(_0044_),
    .CK(clknet_4_11_0_clk),
    .Q(\aso.p[2] ),
    .QN(_3797_));
 DFF_X1 \aso.p[3]$_SDFF_PP0_  (.D(_0045_),
    .CK(clknet_4_12_0_clk),
    .Q(\aso.p[3] ),
    .QN(_3796_));
 DFF_X1 \aso.p[4]$_SDFF_PP0_  (.D(_0046_),
    .CK(clknet_4_13_0_clk),
    .Q(\aso.p[4] ),
    .QN(_3795_));
 DFF_X1 \aso.p[5]$_SDFF_PP0_  (.D(_0047_),
    .CK(clknet_4_13_0_clk),
    .Q(\aso.p[5] ),
    .QN(_3794_));
 DFF_X1 \aso.p[6]$_SDFF_PP0_  (.D(_0048_),
    .CK(clknet_4_15_0_clk),
    .Q(\aso.p[6] ),
    .QN(_3793_));
 DFF_X1 \aso.p[7]$_SDFF_PP0_  (.D(_0049_),
    .CK(clknet_4_14_0_clk),
    .Q(\aso.p[7] ),
    .QN(_3792_));
 DFF_X1 \aso.p[8]$_SDFF_PP0_  (.D(_0050_),
    .CK(clknet_4_14_0_clk),
    .Q(\aso.p[8] ),
    .QN(_3791_));
 DFF_X1 \aso.p[9]$_SDFF_PP0_  (.D(_0051_),
    .CK(clknet_4_15_0_clk),
    .Q(\aso.p[9] ),
    .QN(_3790_));
 DFF_X1 \aso.z0[0]$_SDFF_PP0_  (.D(net14),
    .CK(clknet_4_14_0_clk),
    .Q(\aso.z0[0] ),
    .QN(_3789_));
 DFF_X1 \aso.z0[10]$_SDFF_PP0_  (.D(net6),
    .CK(clknet_4_6_0_clk),
    .Q(\aso.z0[10] ),
    .QN(_0010_));
 DFF_X1 \aso.z0[1]$_SDFF_PP0_  (.D(net98),
    .CK(clknet_4_5_0_clk),
    .Q(\aso.z0[1] ),
    .QN(_3788_));
 DFF_X1 \aso.z0[2]$_SDFF_PP0_  (.D(net4),
    .CK(clknet_4_6_0_clk),
    .Q(\aso.z0[2] ),
    .QN(_3787_));
 DFF_X1 \aso.z0[3]$_SDFF_PP0_  (.D(net12),
    .CK(clknet_4_6_0_clk),
    .Q(\aso.z0[3] ),
    .QN(_0011_));
 DFF_X1 \aso.z0[4]$_SDFF_PP0_  (.D(net112),
    .CK(clknet_4_13_0_clk),
    .Q(\aso.z0[4] ),
    .QN(_3786_));
 DFF_X1 \aso.z0[5]$_SDFF_PP0_  (.D(net10),
    .CK(clknet_4_15_0_clk),
    .Q(\aso.z0[5] ),
    .QN(_3785_));
 DFF_X1 \aso.z0[6]$_SDFF_PP0_  (.D(net8),
    .CK(clknet_4_6_0_clk),
    .Q(\aso.z0[6] ),
    .QN(_0020_));
 DFF_X1 \aso.z0[7]$_SDFF_PP0_  (.D(net100),
    .CK(clknet_4_13_0_clk),
    .Q(\aso.z0[7] ),
    .QN(_3784_));
 DFF_X1 \aso.z0[8]$_SDFF_PP0_  (.D(net104),
    .CK(clknet_4_13_0_clk),
    .Q(\aso.z0[8] ),
    .QN(_3783_));
 DFF_X1 \aso.z0[9]$_SDFF_PP0_  (.D(net2),
    .CK(clknet_4_13_0_clk),
    .Q(\aso.z0[9] ),
    .QN(_3782_));
 DFF_X1 \aso.z1[0]$_SDFF_PP0_  (.D(_0063_),
    .CK(clknet_4_4_0_clk),
    .Q(\aso.z1[0] ),
    .QN(_3781_));
 DFF_X1 \aso.z1[10]$_SDFF_PP0_  (.D(net117),
    .CK(clknet_4_15_0_clk),
    .Q(\aso.z1[10] ),
    .QN(_3780_));
 DFF_X1 \aso.z1[1]$_SDFF_PP0_  (.D(_0065_),
    .CK(clknet_4_7_0_clk),
    .Q(\aso.z1[1] ),
    .QN(_3779_));
 DFF_X1 \aso.z1[2]$_SDFF_PP0_  (.D(_0066_),
    .CK(clknet_4_7_0_clk),
    .Q(\aso.z1[2] ),
    .QN(_3778_));
 DFF_X1 \aso.z1[3]$_SDFF_PP0_  (.D(net125),
    .CK(clknet_4_7_0_clk),
    .Q(\aso.z1[3] ),
    .QN(_3777_));
 DFF_X1 \aso.z1[4]$_SDFF_PP0_  (.D(_0068_),
    .CK(clknet_4_7_0_clk),
    .Q(\aso.z1[4] ),
    .QN(_3776_));
 DFF_X1 \aso.z1[5]$_SDFF_PP0_  (.D(_0069_),
    .CK(clknet_4_5_0_clk),
    .Q(\aso.z1[5] ),
    .QN(_3775_));
 DFF_X1 \aso.z1[6]$_SDFF_PP0_  (.D(_0070_),
    .CK(clknet_4_6_0_clk),
    .Q(\aso.z1[6] ),
    .QN(_3774_));
 DFF_X1 \aso.z1[7]$_SDFF_PP0_  (.D(_0071_),
    .CK(clknet_4_6_0_clk),
    .Q(\aso.z1[7] ),
    .QN(_3773_));
 DFF_X1 \aso.z1[8]$_SDFF_PP0_  (.D(_0072_),
    .CK(clknet_4_15_0_clk),
    .Q(\aso.z1[8] ),
    .QN(_3772_));
 DFF_X1 \aso.z1[9]$_SDFF_PP0_  (.D(_0073_),
    .CK(clknet_4_13_0_clk),
    .Q(\aso.z1[9] ),
    .QN(_3771_));
 DFF_X1 \aso.z2[0]$_SDFF_PP0_  (.D(net74),
    .CK(clknet_4_4_0_clk),
    .Q(\aso.z2[0] ),
    .QN(_3770_));
 DFF_X1 \aso.z2[10]$_SDFF_PP0_  (.D(net62),
    .CK(clknet_4_14_0_clk),
    .Q(\aso.z2[10] ),
    .QN(_3769_));
 DFF_X1 \aso.z2[1]$_SDFF_PP0_  (.D(net44),
    .CK(clknet_4_7_0_clk),
    .Q(\aso.z2[1] ),
    .QN(_3768_));
 DFF_X1 \aso.z2[2]$_SDFF_PP0_  (.D(net40),
    .CK(clknet_4_7_0_clk),
    .Q(\aso.z2[2] ),
    .QN(_3767_));
 DFF_X1 \aso.z2[3]$_SDFF_PP0_  (.D(net60),
    .CK(clknet_4_5_0_clk),
    .Q(\aso.z2[3] ),
    .QN(_3766_));
 DFF_X1 \aso.z2[4]$_SDFF_PP0_  (.D(net34),
    .CK(clknet_4_5_0_clk),
    .Q(\aso.z2[4] ),
    .QN(_3765_));
 DFF_X1 \aso.z2[5]$_SDFF_PP0_  (.D(net28),
    .CK(clknet_4_5_0_clk),
    .Q(\aso.z2[5] ),
    .QN(_3764_));
 DFF_X1 \aso.z2[6]$_SDFF_PP0_  (.D(net22),
    .CK(clknet_4_6_0_clk),
    .Q(\aso.z2[6] ),
    .QN(_3763_));
 DFF_X1 \aso.z2[7]$_SDFF_PP0_  (.D(net24),
    .CK(clknet_4_6_0_clk),
    .Q(\aso.z2[7] ),
    .QN(_3762_));
 DFF_X1 \aso.z2[8]$_SDFF_PP0_  (.D(net66),
    .CK(clknet_4_15_0_clk),
    .Q(\aso.z2[8] ),
    .QN(_3761_));
 DFF_X1 \aso.z2[9]$_SDFF_PP0_  (.D(net36),
    .CK(clknet_4_13_0_clk),
    .Q(\aso.z2[9] ),
    .QN(_3760_));
 DFF_X1 \aso.z3[0]$_SDFF_PP0_  (.D(net58),
    .CK(clknet_4_7_0_clk),
    .Q(\aso.z3[0] ),
    .QN(_3759_));
 DFF_X1 \aso.z3[10]$_SDFF_PP0_  (.D(net48),
    .CK(clknet_4_14_0_clk),
    .Q(\aso.z3[10] ),
    .QN(_3758_));
 DFF_X1 \aso.z3[1]$_SDFF_PP0_  (.D(net26),
    .CK(clknet_4_7_0_clk),
    .Q(\aso.z3[1] ),
    .QN(_3757_));
 DFF_X1 \aso.z3[2]$_SDFF_PP0_  (.D(net54),
    .CK(clknet_4_5_0_clk),
    .Q(\aso.z3[2] ),
    .QN(_3756_));
 DFF_X1 \aso.z3[3]$_SDFF_PP0_  (.D(net46),
    .CK(clknet_4_7_0_clk),
    .Q(\aso.z3[3] ),
    .QN(_3755_));
 DFF_X1 \aso.z3[4]$_SDFF_PP0_  (.D(net32),
    .CK(clknet_4_7_0_clk),
    .Q(\aso.z3[4] ),
    .QN(_3754_));
 DFF_X1 \aso.z3[5]$_SDFF_PP0_  (.D(net18),
    .CK(clknet_4_5_0_clk),
    .Q(\aso.z3[5] ),
    .QN(_3753_));
 DFF_X1 \aso.z3[6]$_SDFF_PP0_  (.D(net20),
    .CK(clknet_4_6_0_clk),
    .Q(\aso.z3[6] ),
    .QN(_3752_));
 DFF_X1 \aso.z3[7]$_SDFF_PP0_  (.D(net42),
    .CK(clknet_4_6_0_clk),
    .Q(\aso.z3[7] ),
    .QN(_3751_));
 DFF_X1 \aso.z3[8]$_SDFF_PP0_  (.D(net30),
    .CK(clknet_4_15_0_clk),
    .Q(\aso.z3[8] ),
    .QN(_3750_));
 DFF_X1 \aso.z3[9]$_SDFF_PP0_  (.D(net38),
    .CK(clknet_4_13_0_clk),
    .Q(\aso.z3[9] ),
    .QN(_3749_));
 DFF_X1 \aso.z4[0]$_SDFF_PP0_  (.D(net68),
    .CK(clknet_4_5_0_clk),
    .Q(\aso.z4[0] ),
    .QN(_3748_));
 DFF_X1 \aso.z4[10]$_SDFF_PP0_  (.D(net90),
    .CK(clknet_4_15_0_clk),
    .Q(\aso.z4[10] ),
    .QN(_3747_));
 DFF_X1 \aso.z4[1]$_SDFF_PP0_  (.D(net80),
    .CK(clknet_4_5_0_clk),
    .Q(\aso.z4[1] ),
    .QN(_3746_));
 DFF_X1 \aso.z4[2]$_SDFF_PP0_  (.D(net92),
    .CK(clknet_4_7_0_clk),
    .Q(\aso.z4[2] ),
    .QN(_3745_));
 DFF_X1 \aso.z4[3]$_SDFF_PP0_  (.D(net86),
    .CK(clknet_4_7_0_clk),
    .Q(\aso.z4[3] ),
    .QN(_3744_));
 DFF_X1 \aso.z4[4]$_SDFF_PP0_  (.D(net84),
    .CK(clknet_4_7_0_clk),
    .Q(\aso.z4[4] ),
    .QN(_3743_));
 DFF_X1 \aso.z4[5]$_SDFF_PP0_  (.D(net72),
    .CK(clknet_4_5_0_clk),
    .Q(\aso.z4[5] ),
    .QN(_3742_));
 DFF_X1 \aso.z4[6]$_SDFF_PP0_  (.D(net50),
    .CK(clknet_4_7_0_clk),
    .Q(\aso.z4[6] ),
    .QN(_3741_));
 DFF_X1 \aso.z4[7]$_SDFF_PP0_  (.D(net78),
    .CK(clknet_4_6_0_clk),
    .Q(\aso.z4[7] ),
    .QN(_3740_));
 DFF_X1 \aso.z4[8]$_SDFF_PP0_  (.D(net56),
    .CK(clknet_4_15_0_clk),
    .Q(\aso.z4[8] ),
    .QN(_3739_));
 DFF_X1 \aso.z4[9]$_SDFF_PP0_  (.D(net16),
    .CK(clknet_4_13_0_clk),
    .Q(\aso.z4[9] ),
    .QN(_3738_));
 DFF_X1 \fir.p0[0]$_SDFF_PP0_  (.D(net110),
    .CK(clknet_4_9_0_clk),
    .Q(\fir.p0[0] ),
    .QN(_3737_));
 DFF_X1 \fir.p0[10]$_SDFF_PP0_  (.D(net94),
    .CK(clknet_4_15_0_clk),
    .Q(\fir.p0[10] ),
    .QN(_3736_));
 DFF_X1 \fir.p0[11]$_SDFF_PP0_  (.D(net96),
    .CK(clknet_4_15_0_clk),
    .Q(\fir.p0[11] ),
    .QN(_3735_));
 DFF_X1 \fir.p0[1]$_SDFF_PP0_  (.D(net52),
    .CK(clknet_4_10_0_clk),
    .Q(\fir.p0[1] ),
    .QN(_3734_));
 DFF_X1 \fir.p0[2]$_SDFF_PP0_  (.D(net70),
    .CK(clknet_4_11_0_clk),
    .Q(\fir.p0[2] ),
    .QN(_3733_));
 DFF_X1 \fir.p0[3]$_SDFF_PP0_  (.D(net88),
    .CK(clknet_4_12_0_clk),
    .Q(\fir.p0[3] ),
    .QN(_3732_));
 DFF_X1 \fir.p0[4]$_SDFF_PP0_  (.D(net106),
    .CK(clknet_4_12_0_clk),
    .Q(\fir.p0[4] ),
    .QN(_3731_));
 DFF_X1 \fir.p0[5]$_SDFF_PP0_  (.D(net108),
    .CK(clknet_4_14_0_clk),
    .Q(\fir.p0[5] ),
    .QN(_3730_));
 DFF_X1 \fir.p0[6]$_SDFF_PP0_  (.D(net76),
    .CK(clknet_4_15_0_clk),
    .Q(\fir.p0[6] ),
    .QN(_3729_));
 DFF_X1 \fir.p0[7]$_SDFF_PP0_  (.D(net82),
    .CK(clknet_4_15_0_clk),
    .Q(\fir.p0[7] ),
    .QN(_3728_));
 DFF_X1 \fir.p0[8]$_SDFF_PP0_  (.D(net64),
    .CK(clknet_4_15_0_clk),
    .Q(\fir.p0[8] ),
    .QN(_3727_));
 DFF_X1 \fir.p0[9]$_SDFF_PP0_  (.D(net102),
    .CK(clknet_4_14_0_clk),
    .Q(\fir.p0[9] ),
    .QN(_0028_));
 DFF_X1 \fir.p1[0]$_SDFF_PP0_  (.D(net154),
    .CK(clknet_4_9_0_clk),
    .Q(\fir.p1[0] ),
    .QN(_0004_));
 DFF_X1 \fir.p1[10]$_SDFF_PP0_  (.D(net156),
    .CK(clknet_4_15_0_clk),
    .Q(\fir.p1[10] ),
    .QN(_3726_));
 DFF_X1 \fir.p1[11]$_SDFF_PP0_  (.D(net130),
    .CK(clknet_4_14_0_clk),
    .Q(\fir.p1[11] ),
    .QN(_0035_));
 DFF_X1 \fir.p1[1]$_SDFF_PP0_  (.D(net162),
    .CK(clknet_4_11_0_clk),
    .Q(\fir.p1[1] ),
    .QN(_0003_));
 DFF_X1 \fir.p1[2]$_SDFF_PP0_  (.D(net178),
    .CK(clknet_4_11_0_clk),
    .Q(\fir.p1[2] ),
    .QN(_0002_));
 DFF_X1 \fir.p1[3]$_SDFF_PP0_  (.D(net204),
    .CK(clknet_4_11_0_clk),
    .Q(\fir.p1[3] ),
    .QN(_0001_));
 DFF_X1 \fir.p1[4]$_SDFF_PP0_  (.D(net234),
    .CK(clknet_4_11_0_clk),
    .Q(\fir.p1[4] ),
    .QN(_0000_));
 DFF_X1 \fir.p1[5]$_SDFF_PP0_  (.D(net208),
    .CK(clknet_4_14_0_clk),
    .Q(\fir.p1[5] ),
    .QN(_0017_));
 DFF_X1 \fir.p1[6]$_SDFF_PP0_  (.D(net236),
    .CK(clknet_4_14_0_clk),
    .Q(\fir.p1[6] ),
    .QN(_0023_));
 DFF_X1 \fir.p1[7]$_SDFF_PP0_  (.D(net226),
    .CK(clknet_4_11_0_clk),
    .Q(\fir.p1[7] ),
    .QN(_3725_));
 DFF_X1 \fir.p1[8]$_SDFF_PP0_  (.D(net228),
    .CK(clknet_4_11_0_clk),
    .Q(\fir.p1[8] ),
    .QN(_3724_));
 DFF_X1 \fir.p1[9]$_SDFF_PP0_  (.D(net127),
    .CK(clknet_4_11_0_clk),
    .Q(\fir.p1[9] ),
    .QN(_3723_));
 DFF_X1 \fir.p2[0]$_SDFF_PP0_  (.D(net114),
    .CK(clknet_4_9_0_clk),
    .Q(\fir.p2[0] ),
    .QN(_0009_));
 DFF_X1 \fir.p2[10]$_SDFF_PP0_  (.D(net206),
    .CK(clknet_4_14_0_clk),
    .Q(\fir.p2[10] ),
    .QN(_3722_));
 DFF_X1 \fir.p2[11]$_SDFF_PP0_  (.D(_0133_),
    .CK(clknet_4_13_0_clk),
    .Q(\fir.p2[11] ),
    .QN(_3721_));
 DFF_X1 \fir.p2[1]$_SDFF_PP0_  (.D(net119),
    .CK(clknet_4_9_0_clk),
    .Q(\fir.p2[1] ),
    .QN(_0008_));
 DFF_X1 \fir.p2[2]$_SDFF_PP0_  (.D(net174),
    .CK(clknet_4_9_0_clk),
    .Q(\fir.p2[2] ),
    .QN(_0007_));
 DFF_X1 \fir.p2[3]$_SDFF_PP0_  (.D(net142),
    .CK(clknet_4_12_0_clk),
    .Q(\fir.p2[3] ),
    .QN(_0006_));
 DFF_X1 \fir.p2[4]$_SDFF_PP0_  (.D(net132),
    .CK(clknet_4_12_0_clk),
    .Q(\fir.p2[4] ),
    .QN(_0019_));
 DFF_X1 \fir.p2[5]$_SDFF_PP0_  (.D(net158),
    .CK(clknet_4_12_0_clk),
    .Q(\fir.p2[5] ),
    .QN(_0025_));
 DFF_X1 \fir.p2[6]$_SDFF_PP0_  (.D(net152),
    .CK(clknet_4_12_0_clk),
    .Q(\fir.p2[6] ),
    .QN(_0005_));
 DFF_X1 \fir.p2[7]$_SDFF_PP0_  (.D(net232),
    .CK(clknet_4_12_0_clk),
    .Q(\fir.p2[7] ),
    .QN(_0018_));
 DFF_X1 \fir.p2[8]$_SDFF_PP0_  (.D(net244),
    .CK(clknet_4_12_0_clk),
    .Q(\fir.p2[8] ),
    .QN(_0024_));
 DFF_X1 \fir.p2[9]$_SDFF_PP0_  (.D(net202),
    .CK(clknet_4_13_0_clk),
    .Q(\fir.p2[9] ),
    .QN(_0038_));
 DFF_X1 \fir.p3[0]$_SDFF_PP0_  (.D(net188),
    .CK(clknet_4_8_0_clk),
    .Q(\fir.p3[0] ),
    .QN(_3720_));
 DFF_X1 \fir.p3[10]$_SDFF_PP0_  (.D(net196),
    .CK(clknet_4_0_0_clk),
    .Q(\fir.p3[10] ),
    .QN(_3719_));
 DFF_X1 \fir.p3[11]$_SDFF_PP0_  (.D(_0145_),
    .CK(clknet_4_4_0_clk),
    .Q(\fir.p3[11] ),
    .QN(_3718_));
 DFF_X1 \fir.p3[1]$_SDFF_PP0_  (.D(net168),
    .CK(clknet_4_8_0_clk),
    .Q(\fir.p3[1] ),
    .QN(_3717_));
 DFF_X1 \fir.p3[2]$_SDFF_PP0_  (.D(net140),
    .CK(clknet_4_9_0_clk),
    .Q(\fir.p3[2] ),
    .QN(_3716_));
 DFF_X1 \fir.p3[3]$_SDFF_PP0_  (.D(net146),
    .CK(clknet_4_9_0_clk),
    .Q(\fir.p3[3] ),
    .QN(_3715_));
 DFF_X1 \fir.p3[4]$_SDFF_PP0_  (.D(net192),
    .CK(clknet_4_3_0_clk),
    .Q(\fir.p3[4] ),
    .QN(_3714_));
 DFF_X1 \fir.p3[5]$_SDFF_PP0_  (.D(net164),
    .CK(clknet_4_3_0_clk),
    .Q(\fir.p3[5] ),
    .QN(_3713_));
 DFF_X1 \fir.p3[6]$_SDFF_PP0_  (.D(net134),
    .CK(clknet_4_3_0_clk),
    .Q(\fir.p3[6] ),
    .QN(_3712_));
 DFF_X1 \fir.p3[7]$_SDFF_PP0_  (.D(net136),
    .CK(clknet_4_4_0_clk),
    .Q(\fir.p3[7] ),
    .QN(_3711_));
 DFF_X1 \fir.p3[8]$_SDFF_PP0_  (.D(net166),
    .CK(clknet_4_6_0_clk),
    .Q(\fir.p3[8] ),
    .QN(_3710_));
 DFF_X1 \fir.p3[9]$_SDFF_PP0_  (.D(net194),
    .CK(clknet_4_3_0_clk),
    .Q(\fir.p3[9] ),
    .QN(_3709_));
 DFF_X1 \fir.p4[0]$_SDFF_PP0_  (.D(net278),
    .CK(clknet_4_8_0_clk),
    .Q(\fir.p4[0] ),
    .QN(_3708_));
 DFF_X1 \fir.p4[10]$_SDFF_PP0_  (.D(net274),
    .CK(clknet_4_4_0_clk),
    .Q(\fir.p4[10] ),
    .QN(_3707_));
 DFF_X1 \fir.p4[11]$_SDFF_PP0_  (.D(_0157_),
    .CK(clknet_4_4_0_clk),
    .Q(\fir.p4[11] ),
    .QN(_0026_));
 DFF_X1 \fir.p4[1]$_SDFF_PP0_  (.D(net270),
    .CK(clknet_4_9_0_clk),
    .Q(\fir.p4[1] ),
    .QN(_3706_));
 DFF_X1 \fir.p4[2]$_SDFF_PP0_  (.D(net210),
    .CK(clknet_4_8_0_clk),
    .Q(\fir.p4[2] ),
    .QN(_3705_));
 DFF_X1 \fir.p4[3]$_SDFF_PP0_  (.D(net248),
    .CK(clknet_4_3_0_clk),
    .Q(\fir.p4[3] ),
    .QN(_3704_));
 DFF_X1 \fir.p4[4]$_SDFF_PP0_  (.D(net212),
    .CK(clknet_4_3_0_clk),
    .Q(\fir.p4[4] ),
    .QN(_3703_));
 DFF_X1 \fir.p4[5]$_SDFF_PP0_  (.D(net246),
    .CK(clknet_4_3_0_clk),
    .Q(\fir.p4[5] ),
    .QN(_3702_));
 DFF_X1 \fir.p4[6]$_SDFF_PP0_  (.D(net218),
    .CK(clknet_4_3_0_clk),
    .Q(\fir.p4[6] ),
    .QN(_3701_));
 DFF_X1 \fir.p4[7]$_SDFF_PP0_  (.D(net222),
    .CK(clknet_4_1_0_clk),
    .Q(\fir.p4[7] ),
    .QN(_3700_));
 DFF_X1 \fir.p4[8]$_SDFF_PP0_  (.D(net220),
    .CK(clknet_4_6_0_clk),
    .Q(\fir.p4[8] ),
    .QN(_3699_));
 DFF_X1 \fir.p4[9]$_SDFF_PP0_  (.D(net272),
    .CK(clknet_4_4_0_clk),
    .Q(\fir.p4[9] ),
    .QN(_3698_));
 DFF_X1 \fir.p5[0]$_SDFF_PP0_  (.D(net276),
    .CK(clknet_4_10_0_clk),
    .Q(\fir.p5[0] ),
    .QN(_0015_));
 DFF_X1 \fir.p5[10]$_SDFF_PP0_  (.D(net242),
    .CK(clknet_4_1_0_clk),
    .Q(\fir.p5[10] ),
    .QN(_3697_));
 DFF_X1 \fir.p5[11]$_SDFF_PP0_  (.D(_0169_),
    .CK(clknet_4_1_0_clk),
    .Q(\fir.p5[11] ),
    .QN(_0029_));
 DFF_X1 \fir.p5[1]$_SDFF_PP0_  (.D(_0170_),
    .CK(clknet_4_8_0_clk),
    .Q(\fir.p5[1] ),
    .QN(_0014_));
 DFF_X1 \fir.p5[2]$_SDFF_PP0_  (.D(net240),
    .CK(clknet_4_8_0_clk),
    .Q(\fir.p5[2] ),
    .QN(_0013_));
 DFF_X1 \fir.p5[3]$_SDFF_PP0_  (.D(net238),
    .CK(clknet_4_2_0_clk),
    .Q(\fir.p5[3] ),
    .QN(_0012_));
 DFF_X1 \fir.p5[4]$_SDFF_PP0_  (.D(net252),
    .CK(clknet_4_2_0_clk),
    .Q(\fir.p5[4] ),
    .QN(_0022_));
 DFF_X1 \fir.p5[5]$_SDFF_PP0_  (.D(net256),
    .CK(clknet_4_0_0_clk),
    .Q(\fir.p5[5] ),
    .QN(_0027_));
 DFF_X1 \fir.p5[6]$_SDFF_PP0_  (.D(net258),
    .CK(clknet_4_0_0_clk),
    .Q(\fir.p5[6] ),
    .QN(_0030_));
 DFF_X1 \fir.p5[7]$_SDFF_PP0_  (.D(net254),
    .CK(clknet_4_1_0_clk),
    .Q(\fir.p5[7] ),
    .QN(_0033_));
 DFF_X1 \fir.p5[8]$_SDFF_PP0_  (.D(_0177_),
    .CK(clknet_4_1_0_clk),
    .Q(\fir.p5[8] ),
    .QN(_0036_));
 DFF_X1 \fir.p5[9]$_SDFF_PP0_  (.D(net262),
    .CK(clknet_4_1_0_clk),
    .Q(\fir.p5[9] ),
    .QN(_0021_));
 DFF_X1 \fir.p6[0]$_SDFF_PP0_  (.D(net184),
    .CK(clknet_4_10_0_clk),
    .Q(\fir.p6[0] ),
    .QN(_3696_));
 DFF_X1 \fir.p6[10]$_SDFF_PP0_  (.D(_0180_),
    .CK(clknet_4_0_0_clk),
    .Q(\fir.p6[10] ),
    .QN(_0039_));
 DFF_X1 \fir.p6[11]$_SDFF_PP0_  (.D(_0181_),
    .CK(clknet_4_1_0_clk),
    .Q(\fir.p6[11] ),
    .QN(_0031_));
 DFF_X1 \fir.p6[1]$_SDFF_PP0_  (.D(net160),
    .CK(clknet_4_10_0_clk),
    .Q(\fir.p6[1] ),
    .QN(_3695_));
 DFF_X1 \fir.p6[2]$_SDFF_PP0_  (.D(net190),
    .CK(clknet_4_10_0_clk),
    .Q(\fir.p6[2] ),
    .QN(_3694_));
 DFF_X1 \fir.p6[3]$_SDFF_PP0_  (.D(net172),
    .CK(clknet_4_10_0_clk),
    .Q(\fir.p6[3] ),
    .QN(_3693_));
 DFF_X1 \fir.p6[4]$_SDFF_PP0_  (.D(net180),
    .CK(clknet_4_10_0_clk),
    .Q(\fir.p6[4] ),
    .QN(_3692_));
 DFF_X1 \fir.p6[5]$_SDFF_PP0_  (.D(net176),
    .CK(clknet_4_8_0_clk),
    .Q(\fir.p6[5] ),
    .QN(_3691_));
 DFF_X1 \fir.p6[6]$_SDFF_PP0_  (.D(_0187_),
    .CK(clknet_4_8_0_clk),
    .Q(\fir.p6[6] ),
    .QN(_3690_));
 DFF_X1 \fir.p6[7]$_SDFF_PP0_  (.D(net198),
    .CK(clknet_4_8_0_clk),
    .Q(\fir.p6[7] ),
    .QN(_0032_));
 DFF_X1 \fir.p6[8]$_SDFF_PP0_  (.D(net182),
    .CK(clknet_4_2_0_clk),
    .Q(\fir.p6[8] ),
    .QN(_0034_));
 DFF_X1 \fir.p6[9]$_SDFF_PP0_  (.D(net200),
    .CK(clknet_4_0_0_clk),
    .Q(\fir.p6[9] ),
    .QN(_0037_));
 DFF_X1 \fir.p7[0]$_SDFF_PP0_  (.D(net122),
    .CK(clknet_4_10_0_clk),
    .Q(\fir.p7[0] ),
    .QN(_3689_));
 DFF_X1 \fir.p7[10]$_SDFF_PP0_  (.D(net138),
    .CK(clknet_4_0_0_clk),
    .Q(\fir.p7[10] ),
    .QN(_3688_));
 DFF_X1 \fir.p7[11]$_SDFF_PP0_  (.D(_0193_),
    .CK(clknet_4_1_0_clk),
    .Q(\fir.p7[11] ),
    .QN(_0016_));
 DFF_X1 \fir.p7[1]$_SDFF_PP0_  (.D(_0194_),
    .CK(clknet_4_10_0_clk),
    .Q(\fir.p7[1] ),
    .QN(_3687_));
 DFF_X1 \fir.p7[2]$_SDFF_PP0_  (.D(net216),
    .CK(clknet_4_10_0_clk),
    .Q(\fir.p7[2] ),
    .QN(_3686_));
 DFF_X1 \fir.p7[3]$_SDFF_PP0_  (.D(net260),
    .CK(clknet_4_10_0_clk),
    .Q(\fir.p7[3] ),
    .QN(_3685_));
 DFF_X1 \fir.p7[4]$_SDFF_PP0_  (.D(net250),
    .CK(clknet_4_10_0_clk),
    .Q(\fir.p7[4] ),
    .QN(_3684_));
 DFF_X1 \fir.p7[5]$_SDFF_PP0_  (.D(net264),
    .CK(clknet_4_10_0_clk),
    .Q(\fir.p7[5] ),
    .QN(_3683_));
 DFF_X1 \fir.p7[6]$_SDFF_PP0_  (.D(net224),
    .CK(clknet_4_10_0_clk),
    .Q(\fir.p7[6] ),
    .QN(_3682_));
 DFF_X1 \fir.p7[7]$_SDFF_PP0_  (.D(net144),
    .CK(clknet_4_8_0_clk),
    .Q(\fir.p7[7] ),
    .QN(_3681_));
 DFF_X1 \fir.p7[8]$_SDFF_PP0_  (.D(net148),
    .CK(clknet_4_2_0_clk),
    .Q(\fir.p7[8] ),
    .QN(_3680_));
 DFF_X1 \fir.p7[9]$_SDFF_PP0_  (.D(net150),
    .CK(clknet_4_2_0_clk),
    .Q(\fir.p7[9] ),
    .QN(_3679_));
 DFF_X1 \q[0]$_SDFF_PP0_  (.D(_0203_),
    .CK(clknet_4_0_0_clk),
    .Q(q[0]),
    .QN(_3678_));
 DFF_X1 \q[10]$_SDFF_PP0_  (.D(_0204_),
    .CK(clknet_4_11_0_clk),
    .Q(q[10]),
    .QN(_3677_));
 DFF_X1 \q[11]$_SDFF_PP0_  (.D(_0205_),
    .CK(clknet_4_5_0_clk),
    .Q(q[11]),
    .QN(_3676_));
 DFF_X1 \q[1]$_SDFF_PP0_  (.D(_0206_),
    .CK(clknet_4_15_0_clk),
    .Q(q[1]),
    .QN(_3675_));
 DFF_X1 \q[2]$_SDFF_PP0_  (.D(_0207_),
    .CK(clknet_4_10_0_clk),
    .Q(q[2]),
    .QN(_3674_));
 DFF_X1 \q[3]$_SDFF_PP0_  (.D(_0208_),
    .CK(clknet_4_2_0_clk),
    .Q(q[3]),
    .QN(_3673_));
 DFF_X1 \q[4]$_SDFF_PP0_  (.D(_0209_),
    .CK(clknet_4_15_0_clk),
    .Q(q[4]),
    .QN(_3672_));
 DFF_X1 \q[5]$_SDFF_PP0_  (.D(_0210_),
    .CK(clknet_4_10_0_clk),
    .Q(q[5]),
    .QN(_3671_));
 DFF_X1 \q[6]$_SDFF_PP0_  (.D(_0211_),
    .CK(clknet_4_0_0_clk),
    .Q(q[6]),
    .QN(_3670_));
 DFF_X1 \q[7]$_SDFF_PP0_  (.D(_0212_),
    .CK(clknet_4_1_0_clk),
    .Q(q[7]),
    .QN(_3669_));
 DFF_X1 \q[8]$_SDFF_PP0_  (.D(_0213_),
    .CK(clknet_4_7_0_clk),
    .Q(q[8]),
    .QN(_3668_));
 DFF_X1 \q[9]$_SDFF_PP0_  (.D(_0214_),
    .CK(clknet_4_1_0_clk),
    .Q(q[9]),
    .QN(_3667_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_117 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_118 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_119 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_120 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_121 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_122 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_123 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_124 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_125 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_126 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_127 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_128 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_129 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_130 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_131 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_132 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_133 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_134 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_135 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_136 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_137 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_138 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_139 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_140 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_141 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_142 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_143 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_144 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_145 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_146 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_147 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_148 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_149 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_150 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_151 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_152 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_153 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_154 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_155 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_156 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_157 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_158 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_159 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_160 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_161 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_162 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_163 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_164 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_165 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_166 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_167 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_168 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_169 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_170 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_171 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_172 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_173 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_174 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_175 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_176 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_177 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_178 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_179 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_180 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_181 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_182 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_183 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_184 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_185 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_186 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_187 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_188 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_189 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_190 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_191 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_192 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_193 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_194 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_195 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_196 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_197 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_198 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_199 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_200 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_201 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_41_202 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_41_203 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_204 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_205 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_43_206 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_43_207 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_208 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_209 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_45_210 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_45_211 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_212 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_213 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_47_214 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_47_215 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_216 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_217 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_49_218 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_49_219 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_220 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_221 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_222 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_223 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_224 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_225 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_53_226 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_53_227 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_228 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_229 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_55_230 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_55_231 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_232 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_233 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_57_234 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_57_235 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_236 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_237 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_238 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_239 ();
 CLKBUF_X1 hold1 (.A(net291),
    .Z(net1));
 CLKBUF_X1 hold2 (.A(_0062_),
    .Z(net2));
 CLKBUF_X1 hold3 (.A(net293),
    .Z(net3));
 CLKBUF_X1 hold4 (.A(_0055_),
    .Z(net4));
 CLKBUF_X1 hold5 (.A(net295),
    .Z(net5));
 CLKBUF_X1 hold6 (.A(_0053_),
    .Z(net6));
 CLKBUF_X1 hold7 (.A(net297),
    .Z(net7));
 CLKBUF_X1 hold8 (.A(_0059_),
    .Z(net8));
 CLKBUF_X1 hold9 (.A(net299),
    .Z(net9));
 CLKBUF_X1 hold10 (.A(_0058_),
    .Z(net10));
 CLKBUF_X1 hold11 (.A(net351),
    .Z(net11));
 CLKBUF_X1 hold12 (.A(_0056_),
    .Z(net12));
 CLKBUF_X1 hold13 (.A(net383),
    .Z(net13));
 CLKBUF_X1 hold14 (.A(_0052_),
    .Z(net14));
 CLKBUF_X1 hold15 (.A(net309),
    .Z(net15));
 CLKBUF_X1 hold16 (.A(_0106_),
    .Z(net16));
 CLKBUF_X1 hold17 (.A(net303),
    .Z(net17));
 CLKBUF_X1 hold18 (.A(_0091_),
    .Z(net18));
 CLKBUF_X1 hold19 (.A(net301),
    .Z(net19));
 CLKBUF_X1 hold20 (.A(_0092_),
    .Z(net20));
 CLKBUF_X1 hold21 (.A(net305),
    .Z(net21));
 CLKBUF_X1 hold22 (.A(_0081_),
    .Z(net22));
 CLKBUF_X1 hold23 (.A(net313),
    .Z(net23));
 CLKBUF_X1 hold24 (.A(_0082_),
    .Z(net24));
 CLKBUF_X1 hold25 (.A(net323),
    .Z(net25));
 CLKBUF_X1 hold26 (.A(_0087_),
    .Z(net26));
 CLKBUF_X1 hold27 (.A(net307),
    .Z(net27));
 CLKBUF_X1 hold28 (.A(_0080_),
    .Z(net28));
 CLKBUF_X1 hold29 (.A(net333),
    .Z(net29));
 CLKBUF_X1 hold30 (.A(_0094_),
    .Z(net30));
 CLKBUF_X1 hold31 (.A(net345),
    .Z(net31));
 CLKBUF_X1 hold32 (.A(_0090_),
    .Z(net32));
 CLKBUF_X1 hold33 (.A(net311),
    .Z(net33));
 CLKBUF_X1 hold34 (.A(_0079_),
    .Z(net34));
 CLKBUF_X1 hold35 (.A(net325),
    .Z(net35));
 CLKBUF_X1 hold36 (.A(_0084_),
    .Z(net36));
 CLKBUF_X1 hold37 (.A(net321),
    .Z(net37));
 CLKBUF_X1 hold38 (.A(_0095_),
    .Z(net38));
 CLKBUF_X1 hold39 (.A(net315),
    .Z(net39));
 CLKBUF_X1 hold40 (.A(_0077_),
    .Z(net40));
 CLKBUF_X1 hold41 (.A(net331),
    .Z(net41));
 CLKBUF_X1 hold42 (.A(_0093_),
    .Z(net42));
 CLKBUF_X1 hold43 (.A(net317),
    .Z(net43));
 CLKBUF_X1 hold44 (.A(_0076_),
    .Z(net44));
 CLKBUF_X1 hold45 (.A(net353),
    .Z(net45));
 CLKBUF_X1 hold46 (.A(_0089_),
    .Z(net46));
 CLKBUF_X1 hold47 (.A(net355),
    .Z(net47));
 CLKBUF_X1 hold48 (.A(_0086_),
    .Z(net48));
 CLKBUF_X1 hold49 (.A(net367),
    .Z(net49));
 CLKBUF_X1 hold50 (.A(_0103_),
    .Z(net50));
 CLKBUF_X1 hold51 (.A(net341),
    .Z(net51));
 CLKBUF_X1 hold52 (.A(_0110_),
    .Z(net52));
 CLKBUF_X1 hold53 (.A(net359),
    .Z(net53));
 CLKBUF_X1 hold54 (.A(_0088_),
    .Z(net54));
 CLKBUF_X1 hold55 (.A(net337),
    .Z(net55));
 CLKBUF_X1 hold56 (.A(_0105_),
    .Z(net56));
 CLKBUF_X1 hold57 (.A(net347),
    .Z(net57));
 CLKBUF_X1 hold58 (.A(_0085_),
    .Z(net58));
 CLKBUF_X1 hold59 (.A(net329),
    .Z(net59));
 CLKBUF_X1 hold60 (.A(_0078_),
    .Z(net60));
 CLKBUF_X1 hold61 (.A(net327),
    .Z(net61));
 CLKBUF_X1 hold62 (.A(_0075_),
    .Z(net62));
 CLKBUF_X1 hold63 (.A(net319),
    .Z(net63));
 CLKBUF_X1 hold64 (.A(_0117_),
    .Z(net64));
 CLKBUF_X1 hold65 (.A(net335),
    .Z(net65));
 CLKBUF_X1 hold66 (.A(_0083_),
    .Z(net66));
 CLKBUF_X1 hold67 (.A(net363),
    .Z(net67));
 CLKBUF_X1 hold68 (.A(_0096_),
    .Z(net68));
 CLKBUF_X1 hold69 (.A(net343),
    .Z(net69));
 CLKBUF_X1 hold70 (.A(_0111_),
    .Z(net70));
 CLKBUF_X1 hold71 (.A(net365),
    .Z(net71));
 CLKBUF_X1 hold72 (.A(_0102_),
    .Z(net72));
 CLKBUF_X1 hold73 (.A(net349),
    .Z(net73));
 CLKBUF_X1 hold74 (.A(_0074_),
    .Z(net74));
 CLKBUF_X1 hold75 (.A(net339),
    .Z(net75));
 CLKBUF_X1 hold76 (.A(_0115_),
    .Z(net76));
 CLKBUF_X1 hold77 (.A(net377),
    .Z(net77));
 CLKBUF_X1 hold78 (.A(_0104_),
    .Z(net78));
 CLKBUF_X1 hold79 (.A(net361),
    .Z(net79));
 CLKBUF_X1 hold80 (.A(_0098_),
    .Z(net80));
 CLKBUF_X1 hold81 (.A(net357),
    .Z(net81));
 CLKBUF_X1 hold82 (.A(_0116_),
    .Z(net82));
 CLKBUF_X1 hold83 (.A(net373),
    .Z(net83));
 CLKBUF_X1 hold84 (.A(_0101_),
    .Z(net84));
 CLKBUF_X1 hold85 (.A(net371),
    .Z(net85));
 CLKBUF_X1 hold86 (.A(_0100_),
    .Z(net86));
 CLKBUF_X1 hold87 (.A(net369),
    .Z(net87));
 CLKBUF_X1 hold88 (.A(_0112_),
    .Z(net88));
 CLKBUF_X1 hold89 (.A(net375),
    .Z(net89));
 CLKBUF_X1 hold90 (.A(_0097_),
    .Z(net90));
 CLKBUF_X1 hold91 (.A(net379),
    .Z(net91));
 CLKBUF_X1 hold92 (.A(_0099_),
    .Z(net92));
 CLKBUF_X1 hold93 (.A(net381),
    .Z(net93));
 CLKBUF_X1 hold94 (.A(_0108_),
    .Z(net94));
 CLKBUF_X1 hold95 (.A(net385),
    .Z(net95));
 CLKBUF_X1 hold96 (.A(_0109_),
    .Z(net96));
 CLKBUF_X1 hold97 (.A(net387),
    .Z(net97));
 CLKBUF_X1 hold98 (.A(_0054_),
    .Z(net98));
 CLKBUF_X1 hold99 (.A(net391),
    .Z(net99));
 CLKBUF_X1 hold100 (.A(_0060_),
    .Z(net100));
 CLKBUF_X1 hold101 (.A(net389),
    .Z(net101));
 CLKBUF_X1 hold102 (.A(_0118_),
    .Z(net102));
 CLKBUF_X1 hold103 (.A(net397),
    .Z(net103));
 CLKBUF_X1 hold104 (.A(_0061_),
    .Z(net104));
 CLKBUF_X1 hold105 (.A(net393),
    .Z(net105));
 CLKBUF_X1 hold106 (.A(_0113_),
    .Z(net106));
 CLKBUF_X1 hold107 (.A(net395),
    .Z(net107));
 CLKBUF_X1 hold108 (.A(_0114_),
    .Z(net108));
 CLKBUF_X1 hold109 (.A(net401),
    .Z(net109));
 CLKBUF_X1 hold110 (.A(_0107_),
    .Z(net110));
 CLKBUF_X1 hold111 (.A(net399),
    .Z(net111));
 CLKBUF_X1 hold112 (.A(_0057_),
    .Z(net112));
 CLKBUF_X1 hold113 (.A(net402),
    .Z(net113));
 CLKBUF_X1 hold114 (.A(_0131_),
    .Z(net114));
 CLKBUF_X1 hold115 (.A(net477),
    .Z(net115));
 CLKBUF_X1 hold116 (.A(_2279_),
    .Z(net116));
 CLKBUF_X1 hold117 (.A(_0064_),
    .Z(net117));
 CLKBUF_X1 hold118 (.A(net403),
    .Z(net118));
 CLKBUF_X1 hold119 (.A(_0134_),
    .Z(net119));
 CLKBUF_X1 hold120 (.A(\fir.p6[0] ),
    .Z(net120));
 CLKBUF_X1 hold121 (.A(_1924_),
    .Z(net121));
 CLKBUF_X1 hold122 (.A(_0191_),
    .Z(net122));
 CLKBUF_X1 hold123 (.A(\aso.z0[3] ),
    .Z(net123));
 CLKBUF_X1 hold124 (.A(_2276_),
    .Z(net124));
 CLKBUF_X1 hold125 (.A(_0067_),
    .Z(net125));
 CLKBUF_X1 hold126 (.A(net409),
    .Z(net126));
 CLKBUF_X1 hold127 (.A(_0130_),
    .Z(net127));
 CLKBUF_X1 hold128 (.A(\fir.p0[11] ),
    .Z(net128));
 CLKBUF_X1 hold129 (.A(_1483_),
    .Z(net129));
 CLKBUF_X1 hold130 (.A(_0121_),
    .Z(net130));
 CLKBUF_X1 hold131 (.A(net404),
    .Z(net131));
 CLKBUF_X1 hold132 (.A(_0137_),
    .Z(net132));
 CLKBUF_X1 hold133 (.A(net420),
    .Z(net133));
 CLKBUF_X1 hold134 (.A(_0151_),
    .Z(net134));
 CLKBUF_X1 hold135 (.A(net417),
    .Z(net135));
 CLKBUF_X1 hold136 (.A(_0152_),
    .Z(net136));
 CLKBUF_X1 hold137 (.A(net405),
    .Z(net137));
 CLKBUF_X1 hold138 (.A(_0192_),
    .Z(net138));
 CLKBUF_X1 hold139 (.A(net411),
    .Z(net139));
 CLKBUF_X1 hold140 (.A(_0147_),
    .Z(net140));
 CLKBUF_X1 hold141 (.A(net421),
    .Z(net141));
 CLKBUF_X1 hold142 (.A(_0136_),
    .Z(net142));
 CLKBUF_X1 hold143 (.A(net406),
    .Z(net143));
 CLKBUF_X1 hold144 (.A(_0200_),
    .Z(net144));
 CLKBUF_X1 hold145 (.A(net416),
    .Z(net145));
 CLKBUF_X1 hold146 (.A(_0148_),
    .Z(net146));
 CLKBUF_X1 hold147 (.A(net407),
    .Z(net147));
 CLKBUF_X1 hold148 (.A(_0201_),
    .Z(net148));
 CLKBUF_X1 hold149 (.A(net408),
    .Z(net149));
 CLKBUF_X1 hold150 (.A(_0202_),
    .Z(net150));
 CLKBUF_X1 hold151 (.A(net414),
    .Z(net151));
 CLKBUF_X1 hold152 (.A(_0139_),
    .Z(net152));
 CLKBUF_X1 hold153 (.A(net413),
    .Z(net153));
 CLKBUF_X1 hold154 (.A(_0119_),
    .Z(net154));
 CLKBUF_X1 hold155 (.A(net412),
    .Z(net155));
 CLKBUF_X1 hold156 (.A(_0120_),
    .Z(net156));
 CLKBUF_X1 hold157 (.A(net415),
    .Z(net157));
 CLKBUF_X1 hold158 (.A(_0138_),
    .Z(net158));
 CLKBUF_X1 hold159 (.A(net425),
    .Z(net159));
 CLKBUF_X1 hold160 (.A(_0182_),
    .Z(net160));
 CLKBUF_X1 hold161 (.A(net410),
    .Z(net161));
 CLKBUF_X1 hold162 (.A(_0122_),
    .Z(net162));
 CLKBUF_X1 hold163 (.A(net422),
    .Z(net163));
 CLKBUF_X1 hold164 (.A(_0150_),
    .Z(net164));
 CLKBUF_X1 hold165 (.A(net424),
    .Z(net165));
 CLKBUF_X1 hold166 (.A(_0153_),
    .Z(net166));
 CLKBUF_X1 hold167 (.A(net418),
    .Z(net167));
 CLKBUF_X1 hold168 (.A(_0146_),
    .Z(net168));
 CLKBUF_X1 hold169 (.A(net439),
    .Z(net169));
 CLKBUF_X1 hold170 (.A(_1536_),
    .Z(net170));
 CLKBUF_X1 hold171 (.A(net427),
    .Z(net171));
 CLKBUF_X1 hold172 (.A(_0184_),
    .Z(net172));
 CLKBUF_X1 hold173 (.A(net423),
    .Z(net173));
 CLKBUF_X1 hold174 (.A(_0135_),
    .Z(net174));
 CLKBUF_X1 hold175 (.A(net434),
    .Z(net175));
 CLKBUF_X1 hold176 (.A(_0186_),
    .Z(net176));
 CLKBUF_X1 hold177 (.A(net419),
    .Z(net177));
 CLKBUF_X1 hold178 (.A(_0123_),
    .Z(net178));
 CLKBUF_X1 hold179 (.A(net428),
    .Z(net179));
 CLKBUF_X1 hold180 (.A(_0185_),
    .Z(net180));
 CLKBUF_X1 hold181 (.A(net432),
    .Z(net181));
 CLKBUF_X1 hold182 (.A(_0189_),
    .Z(net182));
 CLKBUF_X1 hold183 (.A(net435),
    .Z(net183));
 CLKBUF_X1 hold184 (.A(_0179_),
    .Z(net184));
 CLKBUF_X1 hold185 (.A(net454),
    .Z(net185));
 CLKBUF_X1 hold186 (.A(_0705_),
    .Z(net186));
 CLKBUF_X1 hold187 (.A(net446),
    .Z(net187));
 CLKBUF_X1 hold188 (.A(_0143_),
    .Z(net188));
 CLKBUF_X1 hold189 (.A(net433),
    .Z(net189));
 CLKBUF_X1 hold190 (.A(_0183_),
    .Z(net190));
 CLKBUF_X1 hold191 (.A(net426),
    .Z(net191));
 CLKBUF_X1 hold192 (.A(_0149_),
    .Z(net192));
 CLKBUF_X1 hold193 (.A(net451),
    .Z(net193));
 CLKBUF_X1 hold194 (.A(_0154_),
    .Z(net194));
 CLKBUF_X1 hold195 (.A(net455),
    .Z(net195));
 CLKBUF_X1 hold196 (.A(_0144_),
    .Z(net196));
 CLKBUF_X1 hold197 (.A(net431),
    .Z(net197));
 CLKBUF_X1 hold198 (.A(_0188_),
    .Z(net198));
 CLKBUF_X1 hold199 (.A(net429),
    .Z(net199));
 CLKBUF_X1 hold200 (.A(_0190_),
    .Z(net200));
 CLKBUF_X1 hold201 (.A(net437),
    .Z(net201));
 CLKBUF_X1 hold202 (.A(_0142_),
    .Z(net202));
 CLKBUF_X1 hold203 (.A(net442),
    .Z(net203));
 CLKBUF_X1 hold204 (.A(_0124_),
    .Z(net204));
 CLKBUF_X1 hold205 (.A(net443),
    .Z(net205));
 CLKBUF_X1 hold206 (.A(_0132_),
    .Z(net206));
 CLKBUF_X1 hold207 (.A(net436),
    .Z(net207));
 CLKBUF_X1 hold208 (.A(_0126_),
    .Z(net208));
 CLKBUF_X1 hold209 (.A(net440),
    .Z(net209));
 CLKBUF_X1 hold210 (.A(_0159_),
    .Z(net210));
 CLKBUF_X1 hold211 (.A(net438),
    .Z(net211));
 CLKBUF_X1 hold212 (.A(_0161_),
    .Z(net212));
 CLKBUF_X1 hold213 (.A(net470),
    .Z(net213));
 CLKBUF_X1 hold214 (.A(_1904_),
    .Z(net214));
 CLKBUF_X1 hold215 (.A(net441),
    .Z(net215));
 CLKBUF_X1 hold216 (.A(_0195_),
    .Z(net216));
 CLKBUF_X1 hold217 (.A(net445),
    .Z(net217));
 CLKBUF_X1 hold218 (.A(_0163_),
    .Z(net218));
 CLKBUF_X1 hold219 (.A(net450),
    .Z(net219));
 CLKBUF_X1 hold220 (.A(_0165_),
    .Z(net220));
 CLKBUF_X1 hold221 (.A(net448),
    .Z(net221));
 CLKBUF_X1 hold222 (.A(_0164_),
    .Z(net222));
 CLKBUF_X1 hold223 (.A(net447),
    .Z(net223));
 CLKBUF_X1 hold224 (.A(_0199_),
    .Z(net224));
 CLKBUF_X1 hold225 (.A(net475),
    .Z(net225));
 CLKBUF_X1 hold226 (.A(_0128_),
    .Z(net226));
 CLKBUF_X1 hold227 (.A(net480),
    .Z(net227));
 CLKBUF_X1 hold228 (.A(_0129_),
    .Z(net228));
 CLKBUF_X1 hold229 (.A(net458),
    .Z(net229));
 CLKBUF_X1 hold230 (.A(_0434_),
    .Z(net230));
 CLKBUF_X1 hold231 (.A(net456),
    .Z(net231));
 CLKBUF_X1 hold232 (.A(_0140_),
    .Z(net232));
 CLKBUF_X1 hold233 (.A(net453),
    .Z(net233));
 CLKBUF_X1 hold234 (.A(_0125_),
    .Z(net234));
 CLKBUF_X1 hold235 (.A(net457),
    .Z(net235));
 CLKBUF_X1 hold236 (.A(_0127_),
    .Z(net236));
 CLKBUF_X1 hold237 (.A(net461),
    .Z(net237));
 CLKBUF_X1 hold238 (.A(_0172_),
    .Z(net238));
 CLKBUF_X1 hold239 (.A(net464),
    .Z(net239));
 CLKBUF_X1 hold240 (.A(_0171_),
    .Z(net240));
 CLKBUF_X1 hold241 (.A(net469),
    .Z(net241));
 CLKBUF_X1 hold242 (.A(_0168_),
    .Z(net242));
 CLKBUF_X1 hold243 (.A(net466),
    .Z(net243));
 CLKBUF_X1 hold244 (.A(_0141_),
    .Z(net244));
 CLKBUF_X1 hold245 (.A(net452),
    .Z(net245));
 CLKBUF_X1 hold246 (.A(_0162_),
    .Z(net246));
 CLKBUF_X1 hold247 (.A(net460),
    .Z(net247));
 CLKBUF_X1 hold248 (.A(_0160_),
    .Z(net248));
 CLKBUF_X1 hold249 (.A(net465),
    .Z(net249));
 CLKBUF_X1 hold250 (.A(_0197_),
    .Z(net250));
 CLKBUF_X1 hold251 (.A(net463),
    .Z(net251));
 CLKBUF_X1 hold252 (.A(_0173_),
    .Z(net252));
 CLKBUF_X1 hold253 (.A(net467),
    .Z(net253));
 CLKBUF_X1 hold254 (.A(_0176_),
    .Z(net254));
 CLKBUF_X1 hold255 (.A(net471),
    .Z(net255));
 CLKBUF_X1 hold256 (.A(_0174_),
    .Z(net256));
 CLKBUF_X1 hold257 (.A(net472),
    .Z(net257));
 CLKBUF_X1 hold258 (.A(_0175_),
    .Z(net258));
 CLKBUF_X1 hold259 (.A(net473),
    .Z(net259));
 CLKBUF_X1 hold260 (.A(_0196_),
    .Z(net260));
 CLKBUF_X1 hold261 (.A(net479),
    .Z(net261));
 CLKBUF_X1 hold262 (.A(_0178_),
    .Z(net262));
 CLKBUF_X1 hold263 (.A(net462),
    .Z(net263));
 CLKBUF_X1 hold264 (.A(_0198_),
    .Z(net264));
 CLKBUF_X1 hold265 (.A(net486),
    .Z(net265));
 CLKBUF_X1 hold266 (.A(_0921_),
    .Z(net266));
 CLKBUF_X1 hold267 (.A(net484),
    .Z(net267));
 CLKBUF_X1 hold268 (.A(_3517_),
    .Z(net268));
 CLKBUF_X1 hold269 (.A(net468),
    .Z(net269));
 CLKBUF_X1 hold270 (.A(_0158_),
    .Z(net270));
 CLKBUF_X1 hold271 (.A(net474),
    .Z(net271));
 CLKBUF_X1 hold272 (.A(_0166_),
    .Z(net272));
 CLKBUF_X1 hold273 (.A(net483),
    .Z(net273));
 CLKBUF_X1 hold274 (.A(_0156_),
    .Z(net274));
 CLKBUF_X1 hold275 (.A(net487),
    .Z(net275));
 CLKBUF_X1 hold276 (.A(_0167_),
    .Z(net276));
 CLKBUF_X1 hold277 (.A(net488),
    .Z(net277));
 CLKBUF_X1 hold278 (.A(_0155_),
    .Z(net278));
 CLKBUF_X1 hold279 (.A(\fir.p4[1] ),
    .Z(net279));
 CLKBUF_X1 hold280 (.A(_3221_),
    .Z(net280));
 CLKBUF_X1 hold281 (.A(\aso.z0[6] ),
    .Z(net281));
 CLKBUF_X1 hold282 (.A(_2274_),
    .Z(net282));
 CLKBUF_X1 hold283 (.A(net485),
    .Z(net283));
 CLKBUF_X1 hold284 (.A(net478),
    .Z(net284));
 CLKBUF_X1 hold285 (.A(net482),
    .Z(net285));
 CLKBUF_X1 hold286 (.A(net481),
    .Z(net286));
 CLKBUF_X1 hold287 (.A(\aso.z0[0] ),
    .Z(net287));
 CLKBUF_X1 hold288 (.A(\aso.z0[8] ),
    .Z(net288));
 CLKBUF_X1 hold289 (.A(\aso.z0[5] ),
    .Z(net289));
 CLKBUF_X1 hold290 (.A(\aso.z0[9] ),
    .Z(net290));
 CLKBUF_X1 hold291 (.A(z[9]),
    .Z(net291));
 CLKBUF_X1 hold292 (.A(net1),
    .Z(net292));
 CLKBUF_X1 hold293 (.A(z[2]),
    .Z(net293));
 CLKBUF_X1 hold294 (.A(net3),
    .Z(net294));
 CLKBUF_X1 hold295 (.A(z[10]),
    .Z(net295));
 CLKBUF_X1 hold296 (.A(net5),
    .Z(net296));
 CLKBUF_X1 hold297 (.A(z[6]),
    .Z(net297));
 CLKBUF_X1 hold298 (.A(net7),
    .Z(net298));
 CLKBUF_X1 hold299 (.A(z[5]),
    .Z(net299));
 CLKBUF_X1 hold300 (.A(net9),
    .Z(net300));
 CLKBUF_X1 hold301 (.A(\aso.z2[6] ),
    .Z(net301));
 CLKBUF_X1 hold302 (.A(net19),
    .Z(net302));
 CLKBUF_X1 hold303 (.A(\aso.z2[5] ),
    .Z(net303));
 CLKBUF_X1 hold304 (.A(net17),
    .Z(net304));
 CLKBUF_X1 hold305 (.A(\aso.z1[6] ),
    .Z(net305));
 CLKBUF_X1 hold306 (.A(net21),
    .Z(net306));
 CLKBUF_X1 hold307 (.A(\aso.z1[5] ),
    .Z(net307));
 CLKBUF_X1 hold308 (.A(net27),
    .Z(net308));
 CLKBUF_X1 hold309 (.A(\aso.z3[9] ),
    .Z(net309));
 CLKBUF_X1 hold310 (.A(net15),
    .Z(net310));
 CLKBUF_X1 hold311 (.A(\aso.z1[4] ),
    .Z(net311));
 CLKBUF_X1 hold312 (.A(net33),
    .Z(net312));
 CLKBUF_X1 hold313 (.A(\aso.z1[7] ),
    .Z(net313));
 CLKBUF_X1 hold314 (.A(net23),
    .Z(net314));
 CLKBUF_X1 hold315 (.A(\aso.z1[2] ),
    .Z(net315));
 CLKBUF_X1 hold316 (.A(net39),
    .Z(net316));
 CLKBUF_X1 hold317 (.A(\aso.z1[1] ),
    .Z(net317));
 CLKBUF_X1 hold318 (.A(net43),
    .Z(net318));
 CLKBUF_X1 hold319 (.A(\aso.p[8] ),
    .Z(net319));
 CLKBUF_X1 hold320 (.A(net63),
    .Z(net320));
 CLKBUF_X1 hold321 (.A(\aso.z2[9] ),
    .Z(net321));
 CLKBUF_X1 hold322 (.A(net37),
    .Z(net322));
 CLKBUF_X1 hold323 (.A(\aso.z2[1] ),
    .Z(net323));
 CLKBUF_X1 hold324 (.A(net25),
    .Z(net324));
 CLKBUF_X1 hold325 (.A(\aso.z1[9] ),
    .Z(net325));
 CLKBUF_X1 hold326 (.A(net35),
    .Z(net326));
 CLKBUF_X1 hold327 (.A(\aso.z1[10] ),
    .Z(net327));
 CLKBUF_X1 hold328 (.A(net61),
    .Z(net328));
 CLKBUF_X1 hold329 (.A(\aso.z1[3] ),
    .Z(net329));
 CLKBUF_X1 hold330 (.A(net59),
    .Z(net330));
 CLKBUF_X1 hold331 (.A(\aso.z2[7] ),
    .Z(net331));
 CLKBUF_X1 hold332 (.A(net41),
    .Z(net332));
 CLKBUF_X1 hold333 (.A(\aso.z2[8] ),
    .Z(net333));
 CLKBUF_X1 hold334 (.A(net29),
    .Z(net334));
 CLKBUF_X1 hold335 (.A(\aso.z1[8] ),
    .Z(net335));
 CLKBUF_X1 hold336 (.A(net65),
    .Z(net336));
 CLKBUF_X1 hold337 (.A(\aso.z3[8] ),
    .Z(net337));
 CLKBUF_X1 hold338 (.A(net55),
    .Z(net338));
 CLKBUF_X1 hold339 (.A(\aso.p[6] ),
    .Z(net339));
 CLKBUF_X1 hold340 (.A(net75),
    .Z(net340));
 CLKBUF_X1 hold341 (.A(\aso.p[1] ),
    .Z(net341));
 CLKBUF_X1 hold342 (.A(net51),
    .Z(net342));
 CLKBUF_X1 hold343 (.A(\aso.p[2] ),
    .Z(net343));
 CLKBUF_X1 hold344 (.A(net69),
    .Z(net344));
 CLKBUF_X1 hold345 (.A(\aso.z2[4] ),
    .Z(net345));
 CLKBUF_X1 hold346 (.A(net31),
    .Z(net346));
 CLKBUF_X1 hold347 (.A(\aso.z2[0] ),
    .Z(net347));
 CLKBUF_X1 hold348 (.A(net57),
    .Z(net348));
 CLKBUF_X1 hold349 (.A(\aso.z1[0] ),
    .Z(net349));
 CLKBUF_X1 hold350 (.A(net73),
    .Z(net350));
 CLKBUF_X1 hold351 (.A(z[3]),
    .Z(net351));
 CLKBUF_X1 hold352 (.A(net11),
    .Z(net352));
 CLKBUF_X1 hold353 (.A(\aso.z2[3] ),
    .Z(net353));
 CLKBUF_X1 hold354 (.A(net45),
    .Z(net354));
 CLKBUF_X1 hold355 (.A(\aso.z2[10] ),
    .Z(net355));
 CLKBUF_X1 hold356 (.A(net47),
    .Z(net356));
 CLKBUF_X1 hold357 (.A(\aso.p[7] ),
    .Z(net357));
 CLKBUF_X1 hold358 (.A(net81),
    .Z(net358));
 CLKBUF_X1 hold359 (.A(\aso.z2[2] ),
    .Z(net359));
 CLKBUF_X1 hold360 (.A(net53),
    .Z(net360));
 CLKBUF_X1 hold361 (.A(\aso.z3[1] ),
    .Z(net361));
 CLKBUF_X1 hold362 (.A(net79),
    .Z(net362));
 CLKBUF_X1 hold363 (.A(\aso.z3[0] ),
    .Z(net363));
 CLKBUF_X1 hold364 (.A(net67),
    .Z(net364));
 CLKBUF_X1 hold365 (.A(\aso.z3[5] ),
    .Z(net365));
 CLKBUF_X1 hold366 (.A(net71),
    .Z(net366));
 CLKBUF_X1 hold367 (.A(\aso.z3[6] ),
    .Z(net367));
 CLKBUF_X1 hold368 (.A(net49),
    .Z(net368));
 CLKBUF_X1 hold369 (.A(\aso.p[3] ),
    .Z(net369));
 CLKBUF_X1 hold370 (.A(net87),
    .Z(net370));
 CLKBUF_X1 hold371 (.A(\aso.z3[3] ),
    .Z(net371));
 CLKBUF_X1 hold372 (.A(net85),
    .Z(net372));
 CLKBUF_X1 hold373 (.A(\aso.z3[4] ),
    .Z(net373));
 CLKBUF_X1 hold374 (.A(net83),
    .Z(net374));
 CLKBUF_X1 hold375 (.A(\aso.z3[10] ),
    .Z(net375));
 CLKBUF_X1 hold376 (.A(net89),
    .Z(net376));
 CLKBUF_X1 hold377 (.A(\aso.z3[7] ),
    .Z(net377));
 CLKBUF_X1 hold378 (.A(net77),
    .Z(net378));
 CLKBUF_X1 hold379 (.A(\aso.z3[2] ),
    .Z(net379));
 CLKBUF_X1 hold380 (.A(net91),
    .Z(net380));
 CLKBUF_X1 hold381 (.A(\aso.p[10] ),
    .Z(net381));
 CLKBUF_X1 hold382 (.A(net93),
    .Z(net382));
 CLKBUF_X1 hold383 (.A(z[0]),
    .Z(net383));
 CLKBUF_X1 hold384 (.A(net13),
    .Z(net384));
 CLKBUF_X1 hold385 (.A(\aso.p[11] ),
    .Z(net385));
 CLKBUF_X1 hold386 (.A(net95),
    .Z(net386));
 CLKBUF_X1 hold387 (.A(z[1]),
    .Z(net387));
 CLKBUF_X1 hold388 (.A(net97),
    .Z(net388));
 CLKBUF_X1 hold389 (.A(\aso.p[9] ),
    .Z(net389));
 CLKBUF_X1 hold390 (.A(net101),
    .Z(net390));
 CLKBUF_X1 hold391 (.A(z[7]),
    .Z(net391));
 CLKBUF_X1 hold392 (.A(net99),
    .Z(net392));
 CLKBUF_X1 hold393 (.A(\aso.p[4] ),
    .Z(net393));
 CLKBUF_X1 hold394 (.A(net105),
    .Z(net394));
 CLKBUF_X1 hold395 (.A(\aso.p[5] ),
    .Z(net395));
 CLKBUF_X1 hold396 (.A(net107),
    .Z(net396));
 CLKBUF_X1 hold397 (.A(z[8]),
    .Z(net397));
 CLKBUF_X1 hold398 (.A(net103),
    .Z(net398));
 CLKBUF_X1 hold399 (.A(z[4]),
    .Z(net399));
 CLKBUF_X1 hold400 (.A(net111),
    .Z(net400));
 CLKBUF_X1 hold401 (.A(net459),
    .Z(net401));
 CLKBUF_X1 hold402 (.A(net489),
    .Z(net402));
 CLKBUF_X1 hold403 (.A(net476),
    .Z(net403));
 CLKBUF_X1 hold404 (.A(\fir.p1[4] ),
    .Z(net404));
 CLKBUF_X1 hold405 (.A(\fir.p6[10] ),
    .Z(net405));
 CLKBUF_X1 hold406 (.A(\fir.p6[7] ),
    .Z(net406));
 CLKBUF_X1 hold407 (.A(\fir.p6[8] ),
    .Z(net407));
 CLKBUF_X1 hold408 (.A(\fir.p6[9] ),
    .Z(net408));
 CLKBUF_X1 hold409 (.A(\fir.p0[9] ),
    .Z(net409));
 CLKBUF_X1 hold410 (.A(\fir.p0[1] ),
    .Z(net410));
 CLKBUF_X1 hold411 (.A(\fir.p2[2] ),
    .Z(net411));
 CLKBUF_X1 hold412 (.A(\fir.p0[10] ),
    .Z(net412));
 CLKBUF_X1 hold413 (.A(\fir.p0[0] ),
    .Z(net413));
 CLKBUF_X1 hold414 (.A(\fir.p1[6] ),
    .Z(net414));
 CLKBUF_X1 hold415 (.A(\fir.p1[5] ),
    .Z(net415));
 CLKBUF_X1 hold416 (.A(\fir.p2[3] ),
    .Z(net416));
 CLKBUF_X1 hold417 (.A(\fir.p2[7] ),
    .Z(net417));
 CLKBUF_X1 hold418 (.A(\fir.p2[1] ),
    .Z(net418));
 CLKBUF_X1 hold419 (.A(\fir.p0[2] ),
    .Z(net419));
 CLKBUF_X1 hold420 (.A(\fir.p2[6] ),
    .Z(net420));
 BUF_X8 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 BUF_X8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 BUF_X8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 BUF_X8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 BUF_X8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 BUF_X8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 BUF_X8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 BUF_X8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 BUF_X8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 BUF_X8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 BUF_X8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 BUF_X8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 BUF_X8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 BUF_X8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 BUF_X8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 BUF_X8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 BUF_X8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 INV_X8 clkload0 (.A(clknet_4_0_0_clk));
 BUF_X8 clkload1 (.A(clknet_4_1_0_clk));
 INV_X8 clkload2 (.A(clknet_4_2_0_clk));
 INV_X8 clkload3 (.A(clknet_4_3_0_clk));
 INV_X8 clkload4 (.A(clknet_4_4_0_clk));
 BUF_X8 clkload5 (.A(clknet_4_5_0_clk));
 BUF_X4 clkload6 (.A(clknet_4_6_0_clk));
 INV_X2 clkload7 (.A(clknet_4_7_0_clk));
 BUF_X8 clkload8 (.A(clknet_4_8_0_clk));
 INV_X8 clkload9 (.A(clknet_4_9_0_clk));
 BUF_X1 clkload10 (.A(clknet_4_10_0_clk));
 BUF_X8 clkload11 (.A(clknet_4_11_0_clk));
 BUF_X8 clkload12 (.A(clknet_4_12_0_clk));
 INV_X4 clkload13 (.A(clknet_4_13_0_clk));
 INV_X4 clkload14 (.A(clknet_4_14_0_clk));
 CLKBUF_X1 hold421 (.A(\fir.p1[3] ),
    .Z(net421));
 CLKBUF_X1 hold422 (.A(\fir.p2[5] ),
    .Z(net422));
 CLKBUF_X1 hold423 (.A(\fir.p1[2] ),
    .Z(net423));
 CLKBUF_X1 hold424 (.A(\fir.p2[8] ),
    .Z(net424));
 CLKBUF_X1 hold425 (.A(\fir.p5[1] ),
    .Z(net425));
 CLKBUF_X1 hold426 (.A(\fir.p2[4] ),
    .Z(net426));
 CLKBUF_X1 hold427 (.A(\fir.p5[3] ),
    .Z(net427));
 CLKBUF_X1 hold428 (.A(\fir.p5[4] ),
    .Z(net428));
 CLKBUF_X1 hold429 (.A(\fir.p5[9] ),
    .Z(net429));
 CLKBUF_X1 hold430 (.A(\fir.p3[11] ),
    .Z(net430));
 CLKBUF_X1 hold431 (.A(\fir.p5[7] ),
    .Z(net431));
 CLKBUF_X1 hold432 (.A(\fir.p5[8] ),
    .Z(net432));
 CLKBUF_X1 hold433 (.A(\fir.p5[2] ),
    .Z(net433));
 CLKBUF_X1 hold434 (.A(\fir.p5[5] ),
    .Z(net434));
 CLKBUF_X1 hold435 (.A(\fir.p5[0] ),
    .Z(net435));
 CLKBUF_X1 hold436 (.A(\fir.p0[5] ),
    .Z(net436));
 CLKBUF_X1 hold437 (.A(\fir.p1[9] ),
    .Z(net437));
 CLKBUF_X1 hold438 (.A(\fir.p3[4] ),
    .Z(net438));
 CLKBUF_X1 hold439 (.A(\fir.p6[11] ),
    .Z(net439));
 CLKBUF_X1 hold440 (.A(\fir.p3[2] ),
    .Z(net440));
 CLKBUF_X1 hold441 (.A(\fir.p6[2] ),
    .Z(net441));
 CLKBUF_X1 hold442 (.A(\fir.p0[3] ),
    .Z(net442));
 CLKBUF_X1 hold443 (.A(\fir.p1[10] ),
    .Z(net443));
 CLKBUF_X1 hold444 (.A(\fir.p4[11] ),
    .Z(net444));
 CLKBUF_X1 hold445 (.A(\fir.p3[6] ),
    .Z(net445));
 CLKBUF_X1 hold446 (.A(\fir.p2[0] ),
    .Z(net446));
 CLKBUF_X1 hold447 (.A(\fir.p6[6] ),
    .Z(net447));
 CLKBUF_X1 hold448 (.A(\fir.p3[7] ),
    .Z(net448));
 CLKBUF_X1 hold449 (.A(\aso.z0[2] ),
    .Z(net449));
 CLKBUF_X1 hold450 (.A(\fir.p3[8] ),
    .Z(net450));
 CLKBUF_X1 hold451 (.A(\fir.p2[9] ),
    .Z(net451));
 CLKBUF_X1 hold452 (.A(\fir.p3[5] ),
    .Z(net452));
 CLKBUF_X1 hold453 (.A(\fir.p0[4] ),
    .Z(net453));
 CLKBUF_X1 hold454 (.A(\fir.p5[6] ),
    .Z(net454));
 CLKBUF_X1 hold455 (.A(\fir.p2[10] ),
    .Z(net455));
 CLKBUF_X1 hold456 (.A(\fir.p1[7] ),
    .Z(net456));
 CLKBUF_X1 hold457 (.A(\fir.p0[6] ),
    .Z(net457));
 CLKBUF_X1 hold458 (.A(\fir.p5[10] ),
    .Z(net458));
 CLKBUF_X1 hold459 (.A(\aso.p[0] ),
    .Z(net459));
 CLKBUF_X1 hold460 (.A(\fir.p3[3] ),
    .Z(net460));
 CLKBUF_X1 hold461 (.A(\fir.p4[3] ),
    .Z(net461));
 CLKBUF_X1 hold462 (.A(\fir.p6[5] ),
    .Z(net462));
 CLKBUF_X1 hold463 (.A(\fir.p4[4] ),
    .Z(net463));
 CLKBUF_X1 hold464 (.A(\fir.p4[2] ),
    .Z(net464));
 CLKBUF_X1 hold465 (.A(\fir.p6[4] ),
    .Z(net465));
 CLKBUF_X1 hold466 (.A(\fir.p1[8] ),
    .Z(net466));
 CLKBUF_X1 hold467 (.A(\fir.p4[7] ),
    .Z(net467));
 CLKBUF_X1 hold468 (.A(\fir.p3[1] ),
    .Z(net468));
 CLKBUF_X1 hold469 (.A(\fir.p4[10] ),
    .Z(net469));
 CLKBUF_X1 hold470 (.A(\fir.p6[1] ),
    .Z(net470));
 CLKBUF_X1 hold471 (.A(\fir.p4[5] ),
    .Z(net471));
 CLKBUF_X1 hold472 (.A(\fir.p4[6] ),
    .Z(net472));
 CLKBUF_X1 hold473 (.A(\fir.p6[3] ),
    .Z(net473));
 CLKBUF_X1 hold474 (.A(\fir.p3[9] ),
    .Z(net474));
 CLKBUF_X1 hold475 (.A(\fir.p0[7] ),
    .Z(net475));
 CLKBUF_X1 hold476 (.A(\fir.p1[1] ),
    .Z(net476));
 CLKBUF_X1 hold477 (.A(\aso.z0[10] ),
    .Z(net477));
 CLKBUF_X1 hold478 (.A(\aso.z0[7] ),
    .Z(net478));
 CLKBUF_X1 hold479 (.A(\fir.p4[9] ),
    .Z(net479));
 CLKBUF_X1 hold480 (.A(\fir.p0[8] ),
    .Z(net480));
 CLKBUF_X1 hold481 (.A(\fir.p2[11] ),
    .Z(net481));
 CLKBUF_X1 hold482 (.A(\aso.z0[1] ),
    .Z(net482));
 CLKBUF_X1 hold483 (.A(\fir.p3[10] ),
    .Z(net483));
 CLKBUF_X1 hold484 (.A(\fir.p4[8] ),
    .Z(net484));
 CLKBUF_X1 hold485 (.A(\aso.z0[4] ),
    .Z(net485));
 CLKBUF_X1 hold486 (.A(\fir.p1[11] ),
    .Z(net486));
 CLKBUF_X1 hold487 (.A(\fir.p4[0] ),
    .Z(net487));
 CLKBUF_X1 hold488 (.A(\fir.p3[0] ),
    .Z(net488));
 CLKBUF_X1 hold489 (.A(\fir.p1[0] ),
    .Z(net489));
 FILLCELL_X32 FILLER_0_0_1 ();
 FILLCELL_X16 FILLER_0_0_33 ();
 FILLCELL_X1 FILLER_0_0_49 ();
 FILLCELL_X2 FILLER_0_0_57 ();
 FILLCELL_X1 FILLER_0_0_69 ();
 FILLCELL_X8 FILLER_0_0_76 ();
 FILLCELL_X4 FILLER_0_0_84 ();
 FILLCELL_X1 FILLER_0_0_88 ();
 FILLCELL_X4 FILLER_0_0_90 ();
 FILLCELL_X4 FILLER_0_0_107 ();
 FILLCELL_X2 FILLER_0_0_121 ();
 FILLCELL_X1 FILLER_0_0_123 ();
 FILLCELL_X16 FILLER_0_0_127 ();
 FILLCELL_X1 FILLER_0_0_143 ();
 FILLCELL_X2 FILLER_0_0_158 ();
 FILLCELL_X1 FILLER_0_0_160 ();
 FILLCELL_X8 FILLER_0_0_167 ();
 FILLCELL_X2 FILLER_0_0_175 ();
 FILLCELL_X1 FILLER_0_0_177 ();
 FILLCELL_X8 FILLER_0_0_179 ();
 FILLCELL_X4 FILLER_0_0_187 ();
 FILLCELL_X2 FILLER_0_0_191 ();
 FILLCELL_X1 FILLER_0_0_193 ();
 FILLCELL_X2 FILLER_0_0_200 ();
 FILLCELL_X1 FILLER_0_0_202 ();
 FILLCELL_X2 FILLER_0_0_221 ();
 FILLCELL_X1 FILLER_0_0_229 ();
 FILLCELL_X1 FILLER_0_0_233 ();
 FILLCELL_X2 FILLER_0_0_250 ();
 FILLCELL_X2 FILLER_0_0_265 ();
 FILLCELL_X4 FILLER_0_0_271 ();
 FILLCELL_X2 FILLER_0_0_275 ();
 FILLCELL_X1 FILLER_0_0_304 ();
 FILLCELL_X1 FILLER_0_0_311 ();
 FILLCELL_X1 FILLER_0_0_318 ();
 FILLCELL_X1 FILLER_0_0_332 ();
 FILLCELL_X1 FILLER_0_0_336 ();
 FILLCELL_X8 FILLER_0_0_341 ();
 FILLCELL_X4 FILLER_0_0_349 ();
 FILLCELL_X2 FILLER_0_0_353 ();
 FILLCELL_X1 FILLER_0_0_355 ();
 FILLCELL_X32 FILLER_0_0_357 ();
 FILLCELL_X8 FILLER_0_0_389 ();
 FILLCELL_X2 FILLER_0_0_397 ();
 FILLCELL_X4 FILLER_0_0_416 ();
 FILLCELL_X2 FILLER_0_0_420 ();
 FILLCELL_X8 FILLER_0_0_428 ();
 FILLCELL_X4 FILLER_0_0_436 ();
 FILLCELL_X32 FILLER_0_1_1 ();
 FILLCELL_X2 FILLER_0_1_33 ();
 FILLCELL_X1 FILLER_0_1_35 ();
 FILLCELL_X1 FILLER_0_1_46 ();
 FILLCELL_X1 FILLER_0_1_49 ();
 FILLCELL_X1 FILLER_0_1_62 ();
 FILLCELL_X1 FILLER_0_1_73 ();
 FILLCELL_X1 FILLER_0_1_77 ();
 FILLCELL_X2 FILLER_0_1_82 ();
 FILLCELL_X2 FILLER_0_1_90 ();
 FILLCELL_X4 FILLER_0_1_101 ();
 FILLCELL_X1 FILLER_0_1_111 ();
 FILLCELL_X4 FILLER_0_1_118 ();
 FILLCELL_X1 FILLER_0_1_122 ();
 FILLCELL_X1 FILLER_0_1_126 ();
 FILLCELL_X4 FILLER_0_1_133 ();
 FILLCELL_X8 FILLER_0_1_169 ();
 FILLCELL_X1 FILLER_0_1_177 ();
 FILLCELL_X2 FILLER_0_1_185 ();
 FILLCELL_X2 FILLER_0_1_211 ();
 FILLCELL_X2 FILLER_0_1_226 ();
 FILLCELL_X1 FILLER_0_1_228 ();
 FILLCELL_X1 FILLER_0_1_247 ();
 FILLCELL_X4 FILLER_0_1_257 ();
 FILLCELL_X2 FILLER_0_1_271 ();
 FILLCELL_X1 FILLER_0_1_273 ();
 FILLCELL_X2 FILLER_0_1_290 ();
 FILLCELL_X2 FILLER_0_1_295 ();
 FILLCELL_X1 FILLER_0_1_303 ();
 FILLCELL_X2 FILLER_0_1_308 ();
 FILLCELL_X1 FILLER_0_1_310 ();
 FILLCELL_X4 FILLER_0_1_349 ();
 FILLCELL_X2 FILLER_0_1_374 ();
 FILLCELL_X1 FILLER_0_1_379 ();
 FILLCELL_X2 FILLER_0_1_430 ();
 FILLCELL_X4 FILLER_0_1_435 ();
 FILLCELL_X1 FILLER_0_1_439 ();
 FILLCELL_X4 FILLER_0_2_18 ();
 FILLCELL_X2 FILLER_0_2_22 ();
 FILLCELL_X2 FILLER_0_2_47 ();
 FILLCELL_X1 FILLER_0_2_55 ();
 FILLCELL_X2 FILLER_0_2_75 ();
 FILLCELL_X1 FILLER_0_2_83 ();
 FILLCELL_X2 FILLER_0_2_105 ();
 FILLCELL_X2 FILLER_0_2_117 ();
 FILLCELL_X2 FILLER_0_2_153 ();
 FILLCELL_X4 FILLER_0_2_188 ();
 FILLCELL_X2 FILLER_0_2_192 ();
 FILLCELL_X1 FILLER_0_2_200 ();
 FILLCELL_X1 FILLER_0_2_211 ();
 FILLCELL_X8 FILLER_0_2_215 ();
 FILLCELL_X2 FILLER_0_2_223 ();
 FILLCELL_X2 FILLER_0_2_231 ();
 FILLCELL_X1 FILLER_0_2_233 ();
 FILLCELL_X4 FILLER_0_2_238 ();
 FILLCELL_X1 FILLER_0_2_263 ();
 FILLCELL_X1 FILLER_0_2_268 ();
 FILLCELL_X2 FILLER_0_2_271 ();
 FILLCELL_X1 FILLER_0_2_277 ();
 FILLCELL_X4 FILLER_0_2_282 ();
 FILLCELL_X2 FILLER_0_2_286 ();
 FILLCELL_X2 FILLER_0_2_309 ();
 FILLCELL_X1 FILLER_0_2_311 ();
 FILLCELL_X4 FILLER_0_2_318 ();
 FILLCELL_X2 FILLER_0_2_328 ();
 FILLCELL_X2 FILLER_0_2_333 ();
 FILLCELL_X4 FILLER_0_2_338 ();
 FILLCELL_X4 FILLER_0_2_345 ();
 FILLCELL_X8 FILLER_0_2_359 ();
 FILLCELL_X2 FILLER_0_2_421 ();
 FILLCELL_X1 FILLER_0_2_423 ();
 FILLCELL_X16 FILLER_0_3_1 ();
 FILLCELL_X8 FILLER_0_3_17 ();
 FILLCELL_X4 FILLER_0_3_25 ();
 FILLCELL_X8 FILLER_0_3_58 ();
 FILLCELL_X4 FILLER_0_3_66 ();
 FILLCELL_X2 FILLER_0_3_70 ();
 FILLCELL_X1 FILLER_0_3_72 ();
 FILLCELL_X1 FILLER_0_3_78 ();
 FILLCELL_X1 FILLER_0_3_83 ();
 FILLCELL_X1 FILLER_0_3_88 ();
 FILLCELL_X1 FILLER_0_3_95 ();
 FILLCELL_X2 FILLER_0_3_109 ();
 FILLCELL_X1 FILLER_0_3_111 ();
 FILLCELL_X8 FILLER_0_3_115 ();
 FILLCELL_X1 FILLER_0_3_123 ();
 FILLCELL_X16 FILLER_0_3_146 ();
 FILLCELL_X2 FILLER_0_3_162 ();
 FILLCELL_X1 FILLER_0_3_173 ();
 FILLCELL_X1 FILLER_0_3_179 ();
 FILLCELL_X1 FILLER_0_3_184 ();
 FILLCELL_X1 FILLER_0_3_191 ();
 FILLCELL_X1 FILLER_0_3_198 ();
 FILLCELL_X2 FILLER_0_3_205 ();
 FILLCELL_X1 FILLER_0_3_241 ();
 FILLCELL_X2 FILLER_0_3_272 ();
 FILLCELL_X1 FILLER_0_3_286 ();
 FILLCELL_X8 FILLER_0_3_291 ();
 FILLCELL_X2 FILLER_0_3_299 ();
 FILLCELL_X8 FILLER_0_3_310 ();
 FILLCELL_X2 FILLER_0_3_348 ();
 FILLCELL_X1 FILLER_0_3_355 ();
 FILLCELL_X1 FILLER_0_3_369 ();
 FILLCELL_X1 FILLER_0_3_378 ();
 FILLCELL_X2 FILLER_0_3_427 ();
 FILLCELL_X4 FILLER_0_3_436 ();
 FILLCELL_X2 FILLER_0_4_1 ();
 FILLCELL_X1 FILLER_0_4_3 ();
 FILLCELL_X8 FILLER_0_4_12 ();
 FILLCELL_X4 FILLER_0_4_51 ();
 FILLCELL_X2 FILLER_0_4_55 ();
 FILLCELL_X1 FILLER_0_4_64 ();
 FILLCELL_X8 FILLER_0_4_71 ();
 FILLCELL_X2 FILLER_0_4_79 ();
 FILLCELL_X1 FILLER_0_4_81 ();
 FILLCELL_X1 FILLER_0_4_88 ();
 FILLCELL_X2 FILLER_0_4_103 ();
 FILLCELL_X1 FILLER_0_4_105 ();
 FILLCELL_X1 FILLER_0_4_110 ();
 FILLCELL_X4 FILLER_0_4_114 ();
 FILLCELL_X1 FILLER_0_4_118 ();
 FILLCELL_X16 FILLER_0_4_137 ();
 FILLCELL_X4 FILLER_0_4_153 ();
 FILLCELL_X2 FILLER_0_4_157 ();
 FILLCELL_X1 FILLER_0_4_159 ();
 FILLCELL_X8 FILLER_0_4_170 ();
 FILLCELL_X2 FILLER_0_4_178 ();
 FILLCELL_X1 FILLER_0_4_180 ();
 FILLCELL_X4 FILLER_0_4_185 ();
 FILLCELL_X1 FILLER_0_4_195 ();
 FILLCELL_X1 FILLER_0_4_200 ();
 FILLCELL_X1 FILLER_0_4_207 ();
 FILLCELL_X1 FILLER_0_4_211 ();
 FILLCELL_X2 FILLER_0_4_216 ();
 FILLCELL_X8 FILLER_0_4_224 ();
 FILLCELL_X1 FILLER_0_4_232 ();
 FILLCELL_X2 FILLER_0_4_249 ();
 FILLCELL_X8 FILLER_0_4_254 ();
 FILLCELL_X2 FILLER_0_4_262 ();
 FILLCELL_X2 FILLER_0_4_268 ();
 FILLCELL_X16 FILLER_0_4_276 ();
 FILLCELL_X4 FILLER_0_4_298 ();
 FILLCELL_X1 FILLER_0_4_348 ();
 FILLCELL_X2 FILLER_0_4_358 ();
 FILLCELL_X1 FILLER_0_4_390 ();
 FILLCELL_X2 FILLER_0_4_414 ();
 FILLCELL_X1 FILLER_0_4_439 ();
 FILLCELL_X4 FILLER_0_5_1 ();
 FILLCELL_X2 FILLER_0_5_5 ();
 FILLCELL_X1 FILLER_0_5_13 ();
 FILLCELL_X1 FILLER_0_5_18 ();
 FILLCELL_X1 FILLER_0_5_29 ();
 FILLCELL_X1 FILLER_0_5_36 ();
 FILLCELL_X2 FILLER_0_5_43 ();
 FILLCELL_X8 FILLER_0_5_48 ();
 FILLCELL_X1 FILLER_0_5_68 ();
 FILLCELL_X1 FILLER_0_5_72 ();
 FILLCELL_X1 FILLER_0_5_82 ();
 FILLCELL_X2 FILLER_0_5_92 ();
 FILLCELL_X1 FILLER_0_5_109 ();
 FILLCELL_X2 FILLER_0_5_156 ();
 FILLCELL_X1 FILLER_0_5_162 ();
 FILLCELL_X2 FILLER_0_5_197 ();
 FILLCELL_X1 FILLER_0_5_208 ();
 FILLCELL_X1 FILLER_0_5_213 ();
 FILLCELL_X1 FILLER_0_5_220 ();
 FILLCELL_X1 FILLER_0_5_226 ();
 FILLCELL_X4 FILLER_0_5_230 ();
 FILLCELL_X2 FILLER_0_5_234 ();
 FILLCELL_X1 FILLER_0_5_240 ();
 FILLCELL_X4 FILLER_0_5_263 ();
 FILLCELL_X1 FILLER_0_5_267 ();
 FILLCELL_X1 FILLER_0_5_272 ();
 FILLCELL_X2 FILLER_0_5_278 ();
 FILLCELL_X1 FILLER_0_5_280 ();
 FILLCELL_X1 FILLER_0_5_304 ();
 FILLCELL_X2 FILLER_0_5_318 ();
 FILLCELL_X4 FILLER_0_5_343 ();
 FILLCELL_X2 FILLER_0_5_347 ();
 FILLCELL_X4 FILLER_0_5_352 ();
 FILLCELL_X8 FILLER_0_5_411 ();
 FILLCELL_X2 FILLER_0_5_419 ();
 FILLCELL_X1 FILLER_0_5_421 ();
 FILLCELL_X8 FILLER_0_5_429 ();
 FILLCELL_X2 FILLER_0_5_437 ();
 FILLCELL_X1 FILLER_0_5_439 ();
 FILLCELL_X2 FILLER_0_6_1 ();
 FILLCELL_X1 FILLER_0_6_3 ();
 FILLCELL_X1 FILLER_0_6_7 ();
 FILLCELL_X4 FILLER_0_6_27 ();
 FILLCELL_X4 FILLER_0_6_70 ();
 FILLCELL_X1 FILLER_0_6_74 ();
 FILLCELL_X2 FILLER_0_6_81 ();
 FILLCELL_X2 FILLER_0_6_87 ();
 FILLCELL_X1 FILLER_0_6_93 ();
 FILLCELL_X4 FILLER_0_6_98 ();
 FILLCELL_X4 FILLER_0_6_104 ();
 FILLCELL_X2 FILLER_0_6_108 ();
 FILLCELL_X2 FILLER_0_6_130 ();
 FILLCELL_X4 FILLER_0_6_136 ();
 FILLCELL_X1 FILLER_0_6_160 ();
 FILLCELL_X1 FILLER_0_6_167 ();
 FILLCELL_X1 FILLER_0_6_181 ();
 FILLCELL_X2 FILLER_0_6_219 ();
 FILLCELL_X1 FILLER_0_6_253 ();
 FILLCELL_X1 FILLER_0_6_256 ();
 FILLCELL_X1 FILLER_0_6_260 ();
 FILLCELL_X1 FILLER_0_6_274 ();
 FILLCELL_X2 FILLER_0_6_278 ();
 FILLCELL_X1 FILLER_0_6_297 ();
 FILLCELL_X1 FILLER_0_6_301 ();
 FILLCELL_X1 FILLER_0_6_308 ();
 FILLCELL_X1 FILLER_0_6_311 ();
 FILLCELL_X2 FILLER_0_6_318 ();
 FILLCELL_X1 FILLER_0_6_326 ();
 FILLCELL_X1 FILLER_0_6_330 ();
 FILLCELL_X1 FILLER_0_6_334 ();
 FILLCELL_X1 FILLER_0_6_338 ();
 FILLCELL_X1 FILLER_0_6_345 ();
 FILLCELL_X1 FILLER_0_6_366 ();
 FILLCELL_X2 FILLER_0_6_397 ();
 FILLCELL_X8 FILLER_0_7_1 ();
 FILLCELL_X1 FILLER_0_7_9 ();
 FILLCELL_X2 FILLER_0_7_38 ();
 FILLCELL_X4 FILLER_0_7_71 ();
 FILLCELL_X1 FILLER_0_7_75 ();
 FILLCELL_X4 FILLER_0_7_80 ();
 FILLCELL_X1 FILLER_0_7_84 ();
 FILLCELL_X1 FILLER_0_7_107 ();
 FILLCELL_X4 FILLER_0_7_117 ();
 FILLCELL_X8 FILLER_0_7_127 ();
 FILLCELL_X1 FILLER_0_7_135 ();
 FILLCELL_X4 FILLER_0_7_147 ();
 FILLCELL_X1 FILLER_0_7_151 ();
 FILLCELL_X2 FILLER_0_7_158 ();
 FILLCELL_X1 FILLER_0_7_189 ();
 FILLCELL_X4 FILLER_0_7_196 ();
 FILLCELL_X1 FILLER_0_7_200 ();
 FILLCELL_X4 FILLER_0_7_207 ();
 FILLCELL_X1 FILLER_0_7_211 ();
 FILLCELL_X1 FILLER_0_7_215 ();
 FILLCELL_X1 FILLER_0_7_222 ();
 FILLCELL_X2 FILLER_0_7_227 ();
 FILLCELL_X2 FILLER_0_7_239 ();
 FILLCELL_X1 FILLER_0_7_241 ();
 FILLCELL_X1 FILLER_0_7_254 ();
 FILLCELL_X1 FILLER_0_7_289 ();
 FILLCELL_X2 FILLER_0_7_310 ();
 FILLCELL_X8 FILLER_0_7_328 ();
 FILLCELL_X2 FILLER_0_7_340 ();
 FILLCELL_X1 FILLER_0_7_385 ();
 FILLCELL_X1 FILLER_0_7_415 ();
 FILLCELL_X1 FILLER_0_7_436 ();
 FILLCELL_X1 FILLER_0_8_1 ();
 FILLCELL_X1 FILLER_0_8_19 ();
 FILLCELL_X1 FILLER_0_8_24 ();
 FILLCELL_X1 FILLER_0_8_31 ();
 FILLCELL_X1 FILLER_0_8_36 ();
 FILLCELL_X1 FILLER_0_8_43 ();
 FILLCELL_X1 FILLER_0_8_50 ();
 FILLCELL_X8 FILLER_0_8_64 ();
 FILLCELL_X1 FILLER_0_8_72 ();
 FILLCELL_X2 FILLER_0_8_82 ();
 FILLCELL_X1 FILLER_0_8_84 ();
 FILLCELL_X4 FILLER_0_8_115 ();
 FILLCELL_X1 FILLER_0_8_134 ();
 FILLCELL_X2 FILLER_0_8_139 ();
 FILLCELL_X1 FILLER_0_8_141 ();
 FILLCELL_X1 FILLER_0_8_146 ();
 FILLCELL_X1 FILLER_0_8_153 ();
 FILLCELL_X4 FILLER_0_8_179 ();
 FILLCELL_X2 FILLER_0_8_183 ();
 FILLCELL_X2 FILLER_0_8_204 ();
 FILLCELL_X1 FILLER_0_8_206 ();
 FILLCELL_X2 FILLER_0_8_233 ();
 FILLCELL_X2 FILLER_0_8_238 ();
 FILLCELL_X1 FILLER_0_8_240 ();
 FILLCELL_X1 FILLER_0_8_289 ();
 FILLCELL_X1 FILLER_0_8_310 ();
 FILLCELL_X4 FILLER_0_8_321 ();
 FILLCELL_X1 FILLER_0_8_325 ();
 FILLCELL_X1 FILLER_0_8_394 ();
 FILLCELL_X1 FILLER_0_8_398 ();
 FILLCELL_X1 FILLER_0_8_402 ();
 FILLCELL_X1 FILLER_0_8_410 ();
 FILLCELL_X2 FILLER_0_8_438 ();
 FILLCELL_X4 FILLER_0_9_1 ();
 FILLCELL_X2 FILLER_0_9_5 ();
 FILLCELL_X4 FILLER_0_9_22 ();
 FILLCELL_X2 FILLER_0_9_26 ();
 FILLCELL_X4 FILLER_0_9_44 ();
 FILLCELL_X1 FILLER_0_9_48 ();
 FILLCELL_X1 FILLER_0_9_55 ();
 FILLCELL_X1 FILLER_0_9_59 ();
 FILLCELL_X1 FILLER_0_9_66 ();
 FILLCELL_X2 FILLER_0_9_70 ();
 FILLCELL_X2 FILLER_0_9_76 ();
 FILLCELL_X1 FILLER_0_9_91 ();
 FILLCELL_X1 FILLER_0_9_95 ();
 FILLCELL_X2 FILLER_0_9_116 ();
 FILLCELL_X1 FILLER_0_9_118 ();
 FILLCELL_X4 FILLER_0_9_151 ();
 FILLCELL_X2 FILLER_0_9_155 ();
 FILLCELL_X2 FILLER_0_9_160 ();
 FILLCELL_X1 FILLER_0_9_162 ();
 FILLCELL_X2 FILLER_0_9_179 ();
 FILLCELL_X2 FILLER_0_9_185 ();
 FILLCELL_X1 FILLER_0_9_187 ();
 FILLCELL_X2 FILLER_0_9_198 ();
 FILLCELL_X1 FILLER_0_9_200 ();
 FILLCELL_X2 FILLER_0_9_207 ();
 FILLCELL_X2 FILLER_0_9_217 ();
 FILLCELL_X16 FILLER_0_9_233 ();
 FILLCELL_X1 FILLER_0_9_257 ();
 FILLCELL_X2 FILLER_0_9_262 ();
 FILLCELL_X1 FILLER_0_9_270 ();
 FILLCELL_X1 FILLER_0_9_275 ();
 FILLCELL_X1 FILLER_0_9_280 ();
 FILLCELL_X1 FILLER_0_9_284 ();
 FILLCELL_X2 FILLER_0_9_288 ();
 FILLCELL_X1 FILLER_0_9_290 ();
 FILLCELL_X2 FILLER_0_9_294 ();
 FILLCELL_X1 FILLER_0_9_302 ();
 FILLCELL_X1 FILLER_0_9_309 ();
 FILLCELL_X16 FILLER_0_9_320 ();
 FILLCELL_X2 FILLER_0_9_336 ();
 FILLCELL_X2 FILLER_0_9_420 ();
 FILLCELL_X1 FILLER_0_9_426 ();
 FILLCELL_X4 FILLER_0_9_430 ();
 FILLCELL_X1 FILLER_0_10_1 ();
 FILLCELL_X1 FILLER_0_10_8 ();
 FILLCELL_X1 FILLER_0_10_11 ();
 FILLCELL_X1 FILLER_0_10_30 ();
 FILLCELL_X2 FILLER_0_10_39 ();
 FILLCELL_X1 FILLER_0_10_41 ();
 FILLCELL_X2 FILLER_0_10_55 ();
 FILLCELL_X4 FILLER_0_10_60 ();
 FILLCELL_X1 FILLER_0_10_64 ();
 FILLCELL_X1 FILLER_0_10_68 ();
 FILLCELL_X1 FILLER_0_10_74 ();
 FILLCELL_X1 FILLER_0_10_79 ();
 FILLCELL_X1 FILLER_0_10_85 ();
 FILLCELL_X1 FILLER_0_10_101 ();
 FILLCELL_X1 FILLER_0_10_118 ();
 FILLCELL_X2 FILLER_0_10_125 ();
 FILLCELL_X1 FILLER_0_10_127 ();
 FILLCELL_X4 FILLER_0_10_144 ();
 FILLCELL_X2 FILLER_0_10_148 ();
 FILLCELL_X4 FILLER_0_10_177 ();
 FILLCELL_X2 FILLER_0_10_199 ();
 FILLCELL_X1 FILLER_0_10_201 ();
 FILLCELL_X2 FILLER_0_10_205 ();
 FILLCELL_X1 FILLER_0_10_207 ();
 FILLCELL_X2 FILLER_0_10_244 ();
 FILLCELL_X1 FILLER_0_10_246 ();
 FILLCELL_X1 FILLER_0_10_257 ();
 FILLCELL_X1 FILLER_0_10_298 ();
 FILLCELL_X2 FILLER_0_10_307 ();
 FILLCELL_X16 FILLER_0_10_315 ();
 FILLCELL_X1 FILLER_0_10_331 ();
 FILLCELL_X2 FILLER_0_10_344 ();
 FILLCELL_X1 FILLER_0_10_346 ();
 FILLCELL_X1 FILLER_0_10_353 ();
 FILLCELL_X1 FILLER_0_10_362 ();
 FILLCELL_X4 FILLER_0_10_381 ();
 FILLCELL_X1 FILLER_0_10_385 ();
 FILLCELL_X1 FILLER_0_10_395 ();
 FILLCELL_X1 FILLER_0_10_399 ();
 FILLCELL_X1 FILLER_0_10_420 ();
 FILLCELL_X2 FILLER_0_10_438 ();
 FILLCELL_X4 FILLER_0_11_1 ();
 FILLCELL_X2 FILLER_0_11_48 ();
 FILLCELL_X4 FILLER_0_11_73 ();
 FILLCELL_X1 FILLER_0_11_118 ();
 FILLCELL_X4 FILLER_0_11_122 ();
 FILLCELL_X2 FILLER_0_11_126 ();
 FILLCELL_X2 FILLER_0_11_134 ();
 FILLCELL_X1 FILLER_0_11_136 ();
 FILLCELL_X1 FILLER_0_11_140 ();
 FILLCELL_X2 FILLER_0_11_145 ();
 FILLCELL_X1 FILLER_0_11_147 ();
 FILLCELL_X1 FILLER_0_11_158 ();
 FILLCELL_X1 FILLER_0_11_165 ();
 FILLCELL_X2 FILLER_0_11_176 ();
 FILLCELL_X1 FILLER_0_11_179 ();
 FILLCELL_X1 FILLER_0_11_183 ();
 FILLCELL_X1 FILLER_0_11_193 ();
 FILLCELL_X1 FILLER_0_11_221 ();
 FILLCELL_X8 FILLER_0_11_226 ();
 FILLCELL_X1 FILLER_0_11_234 ();
 FILLCELL_X4 FILLER_0_11_238 ();
 FILLCELL_X2 FILLER_0_11_244 ();
 FILLCELL_X4 FILLER_0_11_275 ();
 FILLCELL_X1 FILLER_0_11_279 ();
 FILLCELL_X2 FILLER_0_11_292 ();
 FILLCELL_X1 FILLER_0_11_300 ();
 FILLCELL_X2 FILLER_0_11_315 ();
 FILLCELL_X1 FILLER_0_11_317 ();
 FILLCELL_X2 FILLER_0_11_334 ();
 FILLCELL_X1 FILLER_0_11_341 ();
 FILLCELL_X4 FILLER_0_11_348 ();
 FILLCELL_X1 FILLER_0_11_355 ();
 FILLCELL_X2 FILLER_0_11_387 ();
 FILLCELL_X1 FILLER_0_11_389 ();
 FILLCELL_X1 FILLER_0_11_405 ();
 FILLCELL_X1 FILLER_0_12_1 ();
 FILLCELL_X4 FILLER_0_12_27 ();
 FILLCELL_X1 FILLER_0_12_31 ();
 FILLCELL_X4 FILLER_0_12_41 ();
 FILLCELL_X1 FILLER_0_12_45 ();
 FILLCELL_X1 FILLER_0_12_59 ();
 FILLCELL_X8 FILLER_0_12_63 ();
 FILLCELL_X4 FILLER_0_12_71 ();
 FILLCELL_X2 FILLER_0_12_75 ();
 FILLCELL_X1 FILLER_0_12_84 ();
 FILLCELL_X1 FILLER_0_12_90 ();
 FILLCELL_X1 FILLER_0_12_97 ();
 FILLCELL_X1 FILLER_0_12_106 ();
 FILLCELL_X1 FILLER_0_12_117 ();
 FILLCELL_X1 FILLER_0_12_122 ();
 FILLCELL_X1 FILLER_0_12_128 ();
 FILLCELL_X1 FILLER_0_12_147 ();
 FILLCELL_X1 FILLER_0_12_173 ();
 FILLCELL_X2 FILLER_0_12_180 ();
 FILLCELL_X4 FILLER_0_12_186 ();
 FILLCELL_X2 FILLER_0_12_190 ();
 FILLCELL_X1 FILLER_0_12_192 ();
 FILLCELL_X1 FILLER_0_12_210 ();
 FILLCELL_X1 FILLER_0_12_223 ();
 FILLCELL_X1 FILLER_0_12_230 ();
 FILLCELL_X1 FILLER_0_12_237 ();
 FILLCELL_X2 FILLER_0_12_248 ();
 FILLCELL_X1 FILLER_0_12_250 ();
 FILLCELL_X2 FILLER_0_12_281 ();
 FILLCELL_X1 FILLER_0_12_285 ();
 FILLCELL_X1 FILLER_0_12_292 ();
 FILLCELL_X2 FILLER_0_12_299 ();
 FILLCELL_X1 FILLER_0_12_327 ();
 FILLCELL_X1 FILLER_0_12_330 ();
 FILLCELL_X1 FILLER_0_12_349 ();
 FILLCELL_X1 FILLER_0_12_355 ();
 FILLCELL_X1 FILLER_0_12_380 ();
 FILLCELL_X1 FILLER_0_12_385 ();
 FILLCELL_X1 FILLER_0_12_405 ();
 FILLCELL_X1 FILLER_0_12_426 ();
 FILLCELL_X4 FILLER_0_12_430 ();
 FILLCELL_X2 FILLER_0_12_434 ();
 FILLCELL_X2 FILLER_0_13_25 ();
 FILLCELL_X1 FILLER_0_13_42 ();
 FILLCELL_X2 FILLER_0_13_58 ();
 FILLCELL_X1 FILLER_0_13_60 ();
 FILLCELL_X2 FILLER_0_13_73 ();
 FILLCELL_X1 FILLER_0_13_75 ();
 FILLCELL_X1 FILLER_0_13_84 ();
 FILLCELL_X1 FILLER_0_13_118 ();
 FILLCELL_X2 FILLER_0_13_128 ();
 FILLCELL_X1 FILLER_0_13_141 ();
 FILLCELL_X1 FILLER_0_13_155 ();
 FILLCELL_X2 FILLER_0_13_159 ();
 FILLCELL_X1 FILLER_0_13_161 ();
 FILLCELL_X1 FILLER_0_13_165 ();
 FILLCELL_X4 FILLER_0_13_171 ();
 FILLCELL_X2 FILLER_0_13_175 ();
 FILLCELL_X1 FILLER_0_13_177 ();
 FILLCELL_X4 FILLER_0_13_198 ();
 FILLCELL_X1 FILLER_0_13_216 ();
 FILLCELL_X8 FILLER_0_13_219 ();
 FILLCELL_X4 FILLER_0_13_227 ();
 FILLCELL_X1 FILLER_0_13_231 ();
 FILLCELL_X8 FILLER_0_13_253 ();
 FILLCELL_X2 FILLER_0_13_261 ();
 FILLCELL_X1 FILLER_0_13_272 ();
 FILLCELL_X1 FILLER_0_13_277 ();
 FILLCELL_X1 FILLER_0_13_287 ();
 FILLCELL_X8 FILLER_0_13_298 ();
 FILLCELL_X4 FILLER_0_13_306 ();
 FILLCELL_X2 FILLER_0_13_310 ();
 FILLCELL_X1 FILLER_0_13_321 ();
 FILLCELL_X1 FILLER_0_13_326 ();
 FILLCELL_X1 FILLER_0_13_357 ();
 FILLCELL_X1 FILLER_0_13_413 ();
 FILLCELL_X2 FILLER_0_13_420 ();
 FILLCELL_X1 FILLER_0_13_422 ();
 FILLCELL_X4 FILLER_0_14_1 ();
 FILLCELL_X2 FILLER_0_14_5 ();
 FILLCELL_X1 FILLER_0_14_7 ();
 FILLCELL_X8 FILLER_0_14_17 ();
 FILLCELL_X2 FILLER_0_14_52 ();
 FILLCELL_X4 FILLER_0_14_57 ();
 FILLCELL_X2 FILLER_0_14_61 ();
 FILLCELL_X1 FILLER_0_14_63 ();
 FILLCELL_X1 FILLER_0_14_77 ();
 FILLCELL_X1 FILLER_0_14_81 ();
 FILLCELL_X1 FILLER_0_14_88 ();
 FILLCELL_X2 FILLER_0_14_112 ();
 FILLCELL_X8 FILLER_0_14_120 ();
 FILLCELL_X1 FILLER_0_14_128 ();
 FILLCELL_X4 FILLER_0_14_136 ();
 FILLCELL_X2 FILLER_0_14_140 ();
 FILLCELL_X1 FILLER_0_14_142 ();
 FILLCELL_X1 FILLER_0_14_165 ();
 FILLCELL_X2 FILLER_0_14_187 ();
 FILLCELL_X1 FILLER_0_14_199 ();
 FILLCELL_X4 FILLER_0_14_209 ();
 FILLCELL_X2 FILLER_0_14_232 ();
 FILLCELL_X1 FILLER_0_14_242 ();
 FILLCELL_X4 FILLER_0_14_247 ();
 FILLCELL_X2 FILLER_0_14_251 ();
 FILLCELL_X1 FILLER_0_14_253 ();
 FILLCELL_X4 FILLER_0_14_263 ();
 FILLCELL_X1 FILLER_0_14_290 ();
 FILLCELL_X16 FILLER_0_14_294 ();
 FILLCELL_X2 FILLER_0_14_310 ();
 FILLCELL_X1 FILLER_0_14_312 ();
 FILLCELL_X2 FILLER_0_14_328 ();
 FILLCELL_X1 FILLER_0_14_330 ();
 FILLCELL_X1 FILLER_0_14_337 ();
 FILLCELL_X2 FILLER_0_14_360 ();
 FILLCELL_X1 FILLER_0_14_362 ();
 FILLCELL_X1 FILLER_0_14_368 ();
 FILLCELL_X1 FILLER_0_14_386 ();
 FILLCELL_X8 FILLER_0_14_429 ();
 FILLCELL_X2 FILLER_0_14_437 ();
 FILLCELL_X1 FILLER_0_14_439 ();
 FILLCELL_X1 FILLER_0_15_7 ();
 FILLCELL_X8 FILLER_0_15_12 ();
 FILLCELL_X4 FILLER_0_15_37 ();
 FILLCELL_X2 FILLER_0_15_41 ();
 FILLCELL_X4 FILLER_0_15_46 ();
 FILLCELL_X1 FILLER_0_15_50 ();
 FILLCELL_X2 FILLER_0_15_57 ();
 FILLCELL_X2 FILLER_0_15_62 ();
 FILLCELL_X1 FILLER_0_15_79 ();
 FILLCELL_X1 FILLER_0_15_84 ();
 FILLCELL_X2 FILLER_0_15_106 ();
 FILLCELL_X1 FILLER_0_15_108 ();
 FILLCELL_X8 FILLER_0_15_121 ();
 FILLCELL_X2 FILLER_0_15_129 ();
 FILLCELL_X1 FILLER_0_15_131 ();
 FILLCELL_X1 FILLER_0_15_138 ();
 FILLCELL_X4 FILLER_0_15_142 ();
 FILLCELL_X1 FILLER_0_15_146 ();
 FILLCELL_X1 FILLER_0_15_151 ();
 FILLCELL_X2 FILLER_0_15_158 ();
 FILLCELL_X1 FILLER_0_15_179 ();
 FILLCELL_X1 FILLER_0_15_186 ();
 FILLCELL_X1 FILLER_0_15_189 ();
 FILLCELL_X1 FILLER_0_15_193 ();
 FILLCELL_X1 FILLER_0_15_197 ();
 FILLCELL_X4 FILLER_0_15_214 ();
 FILLCELL_X1 FILLER_0_15_218 ();
 FILLCELL_X2 FILLER_0_15_261 ();
 FILLCELL_X4 FILLER_0_15_271 ();
 FILLCELL_X8 FILLER_0_15_290 ();
 FILLCELL_X4 FILLER_0_15_301 ();
 FILLCELL_X2 FILLER_0_15_305 ();
 FILLCELL_X1 FILLER_0_15_307 ();
 FILLCELL_X2 FILLER_0_15_321 ();
 FILLCELL_X1 FILLER_0_15_323 ();
 FILLCELL_X1 FILLER_0_15_328 ();
 FILLCELL_X1 FILLER_0_15_334 ();
 FILLCELL_X2 FILLER_0_15_339 ();
 FILLCELL_X2 FILLER_0_15_347 ();
 FILLCELL_X4 FILLER_0_15_352 ();
 FILLCELL_X1 FILLER_0_15_390 ();
 FILLCELL_X1 FILLER_0_15_397 ();
 FILLCELL_X4 FILLER_0_16_1 ();
 FILLCELL_X1 FILLER_0_16_22 ();
 FILLCELL_X2 FILLER_0_16_25 ();
 FILLCELL_X1 FILLER_0_16_27 ();
 FILLCELL_X1 FILLER_0_16_38 ();
 FILLCELL_X1 FILLER_0_16_72 ();
 FILLCELL_X2 FILLER_0_16_77 ();
 FILLCELL_X4 FILLER_0_16_85 ();
 FILLCELL_X2 FILLER_0_16_96 ();
 FILLCELL_X2 FILLER_0_16_142 ();
 FILLCELL_X1 FILLER_0_16_144 ();
 FILLCELL_X1 FILLER_0_16_148 ();
 FILLCELL_X2 FILLER_0_16_172 ();
 FILLCELL_X1 FILLER_0_16_177 ();
 FILLCELL_X2 FILLER_0_16_188 ();
 FILLCELL_X4 FILLER_0_16_196 ();
 FILLCELL_X1 FILLER_0_16_210 ();
 FILLCELL_X1 FILLER_0_16_217 ();
 FILLCELL_X1 FILLER_0_16_224 ();
 FILLCELL_X1 FILLER_0_16_235 ();
 FILLCELL_X1 FILLER_0_16_239 ();
 FILLCELL_X1 FILLER_0_16_249 ();
 FILLCELL_X2 FILLER_0_16_284 ();
 FILLCELL_X2 FILLER_0_16_289 ();
 FILLCELL_X1 FILLER_0_16_291 ();
 FILLCELL_X2 FILLER_0_16_315 ();
 FILLCELL_X2 FILLER_0_16_329 ();
 FILLCELL_X1 FILLER_0_16_331 ();
 FILLCELL_X1 FILLER_0_16_362 ();
 FILLCELL_X8 FILLER_0_17_24 ();
 FILLCELL_X1 FILLER_0_17_35 ();
 FILLCELL_X1 FILLER_0_17_50 ();
 FILLCELL_X1 FILLER_0_17_54 ();
 FILLCELL_X2 FILLER_0_17_61 ();
 FILLCELL_X2 FILLER_0_17_69 ();
 FILLCELL_X4 FILLER_0_17_88 ();
 FILLCELL_X1 FILLER_0_17_92 ();
 FILLCELL_X4 FILLER_0_17_96 ();
 FILLCELL_X4 FILLER_0_17_106 ();
 FILLCELL_X2 FILLER_0_17_127 ();
 FILLCELL_X1 FILLER_0_17_132 ();
 FILLCELL_X1 FILLER_0_17_139 ();
 FILLCELL_X2 FILLER_0_17_152 ();
 FILLCELL_X2 FILLER_0_17_176 ();
 FILLCELL_X8 FILLER_0_17_197 ();
 FILLCELL_X4 FILLER_0_17_208 ();
 FILLCELL_X1 FILLER_0_17_212 ();
 FILLCELL_X4 FILLER_0_17_219 ();
 FILLCELL_X2 FILLER_0_17_223 ();
 FILLCELL_X1 FILLER_0_17_225 ();
 FILLCELL_X8 FILLER_0_17_228 ();
 FILLCELL_X1 FILLER_0_17_236 ();
 FILLCELL_X4 FILLER_0_17_243 ();
 FILLCELL_X1 FILLER_0_17_247 ();
 FILLCELL_X4 FILLER_0_17_281 ();
 FILLCELL_X1 FILLER_0_17_289 ();
 FILLCELL_X1 FILLER_0_17_296 ();
 FILLCELL_X2 FILLER_0_17_300 ();
 FILLCELL_X1 FILLER_0_17_306 ();
 FILLCELL_X4 FILLER_0_17_310 ();
 FILLCELL_X1 FILLER_0_17_314 ();
 FILLCELL_X2 FILLER_0_17_327 ();
 FILLCELL_X2 FILLER_0_17_354 ();
 FILLCELL_X1 FILLER_0_17_402 ();
 FILLCELL_X1 FILLER_0_17_409 ();
 FILLCELL_X4 FILLER_0_17_424 ();
 FILLCELL_X1 FILLER_0_17_431 ();
 FILLCELL_X1 FILLER_0_17_439 ();
 FILLCELL_X8 FILLER_0_18_1 ();
 FILLCELL_X4 FILLER_0_18_9 ();
 FILLCELL_X8 FILLER_0_18_59 ();
 FILLCELL_X4 FILLER_0_18_67 ();
 FILLCELL_X1 FILLER_0_18_75 ();
 FILLCELL_X4 FILLER_0_18_83 ();
 FILLCELL_X2 FILLER_0_18_87 ();
 FILLCELL_X16 FILLER_0_18_99 ();
 FILLCELL_X1 FILLER_0_18_127 ();
 FILLCELL_X4 FILLER_0_18_131 ();
 FILLCELL_X1 FILLER_0_18_141 ();
 FILLCELL_X2 FILLER_0_18_155 ();
 FILLCELL_X4 FILLER_0_18_163 ();
 FILLCELL_X2 FILLER_0_18_167 ();
 FILLCELL_X8 FILLER_0_18_176 ();
 FILLCELL_X1 FILLER_0_18_187 ();
 FILLCELL_X1 FILLER_0_18_194 ();
 FILLCELL_X2 FILLER_0_18_220 ();
 FILLCELL_X1 FILLER_0_18_232 ();
 FILLCELL_X1 FILLER_0_18_235 ();
 FILLCELL_X1 FILLER_0_18_240 ();
 FILLCELL_X1 FILLER_0_18_244 ();
 FILLCELL_X1 FILLER_0_18_247 ();
 FILLCELL_X2 FILLER_0_18_252 ();
 FILLCELL_X2 FILLER_0_18_288 ();
 FILLCELL_X4 FILLER_0_18_300 ();
 FILLCELL_X2 FILLER_0_18_304 ();
 FILLCELL_X1 FILLER_0_18_306 ();
 FILLCELL_X2 FILLER_0_18_327 ();
 FILLCELL_X2 FILLER_0_18_366 ();
 FILLCELL_X2 FILLER_0_18_399 ();
 FILLCELL_X1 FILLER_0_18_401 ();
 FILLCELL_X2 FILLER_0_18_431 ();
 FILLCELL_X1 FILLER_0_18_439 ();
 FILLCELL_X8 FILLER_0_19_1 ();
 FILLCELL_X2 FILLER_0_19_9 ();
 FILLCELL_X1 FILLER_0_19_11 ();
 FILLCELL_X2 FILLER_0_19_35 ();
 FILLCELL_X1 FILLER_0_19_37 ();
 FILLCELL_X1 FILLER_0_19_51 ();
 FILLCELL_X8 FILLER_0_19_56 ();
 FILLCELL_X2 FILLER_0_19_64 ();
 FILLCELL_X1 FILLER_0_19_66 ();
 FILLCELL_X1 FILLER_0_19_82 ();
 FILLCELL_X1 FILLER_0_19_107 ();
 FILLCELL_X1 FILLER_0_19_142 ();
 FILLCELL_X2 FILLER_0_19_159 ();
 FILLCELL_X1 FILLER_0_19_161 ();
 FILLCELL_X2 FILLER_0_19_197 ();
 FILLCELL_X1 FILLER_0_19_202 ();
 FILLCELL_X2 FILLER_0_19_206 ();
 FILLCELL_X2 FILLER_0_19_219 ();
 FILLCELL_X1 FILLER_0_19_224 ();
 FILLCELL_X4 FILLER_0_19_229 ();
 FILLCELL_X1 FILLER_0_19_281 ();
 FILLCELL_X4 FILLER_0_19_288 ();
 FILLCELL_X4 FILLER_0_19_298 ();
 FILLCELL_X2 FILLER_0_19_302 ();
 FILLCELL_X2 FILLER_0_19_349 ();
 FILLCELL_X1 FILLER_0_19_351 ();
 FILLCELL_X1 FILLER_0_19_387 ();
 FILLCELL_X1 FILLER_0_19_395 ();
 FILLCELL_X1 FILLER_0_19_413 ();
 FILLCELL_X1 FILLER_0_19_431 ();
 FILLCELL_X4 FILLER_0_19_435 ();
 FILLCELL_X1 FILLER_0_19_439 ();
 FILLCELL_X2 FILLER_0_20_1 ();
 FILLCELL_X1 FILLER_0_20_3 ();
 FILLCELL_X2 FILLER_0_20_28 ();
 FILLCELL_X1 FILLER_0_20_30 ();
 FILLCELL_X4 FILLER_0_20_84 ();
 FILLCELL_X1 FILLER_0_20_88 ();
 FILLCELL_X2 FILLER_0_20_90 ();
 FILLCELL_X2 FILLER_0_20_102 ();
 FILLCELL_X1 FILLER_0_20_104 ();
 FILLCELL_X1 FILLER_0_20_111 ();
 FILLCELL_X1 FILLER_0_20_115 ();
 FILLCELL_X2 FILLER_0_20_129 ();
 FILLCELL_X4 FILLER_0_20_154 ();
 FILLCELL_X4 FILLER_0_20_162 ();
 FILLCELL_X1 FILLER_0_20_166 ();
 FILLCELL_X1 FILLER_0_20_185 ();
 FILLCELL_X1 FILLER_0_20_197 ();
 FILLCELL_X1 FILLER_0_20_201 ();
 FILLCELL_X1 FILLER_0_20_208 ();
 FILLCELL_X1 FILLER_0_20_218 ();
 FILLCELL_X2 FILLER_0_20_222 ();
 FILLCELL_X4 FILLER_0_20_236 ();
 FILLCELL_X1 FILLER_0_20_240 ();
 FILLCELL_X1 FILLER_0_20_245 ();
 FILLCELL_X4 FILLER_0_20_250 ();
 FILLCELL_X8 FILLER_0_20_257 ();
 FILLCELL_X2 FILLER_0_20_265 ();
 FILLCELL_X2 FILLER_0_20_285 ();
 FILLCELL_X1 FILLER_0_20_287 ();
 FILLCELL_X1 FILLER_0_20_296 ();
 FILLCELL_X1 FILLER_0_20_303 ();
 FILLCELL_X1 FILLER_0_20_311 ();
 FILLCELL_X1 FILLER_0_20_318 ();
 FILLCELL_X2 FILLER_0_20_352 ();
 FILLCELL_X1 FILLER_0_20_358 ();
 FILLCELL_X2 FILLER_0_20_421 ();
 FILLCELL_X4 FILLER_0_21_1 ();
 FILLCELL_X2 FILLER_0_21_5 ();
 FILLCELL_X1 FILLER_0_21_7 ();
 FILLCELL_X2 FILLER_0_21_48 ();
 FILLCELL_X4 FILLER_0_21_53 ();
 FILLCELL_X2 FILLER_0_21_57 ();
 FILLCELL_X2 FILLER_0_21_65 ();
 FILLCELL_X8 FILLER_0_21_99 ();
 FILLCELL_X4 FILLER_0_21_107 ();
 FILLCELL_X1 FILLER_0_21_111 ();
 FILLCELL_X2 FILLER_0_21_136 ();
 FILLCELL_X4 FILLER_0_21_188 ();
 FILLCELL_X2 FILLER_0_21_198 ();
 FILLCELL_X2 FILLER_0_21_210 ();
 FILLCELL_X1 FILLER_0_21_212 ();
 FILLCELL_X1 FILLER_0_21_243 ();
 FILLCELL_X2 FILLER_0_21_250 ();
 FILLCELL_X1 FILLER_0_21_252 ();
 FILLCELL_X1 FILLER_0_21_259 ();
 FILLCELL_X4 FILLER_0_21_273 ();
 FILLCELL_X4 FILLER_0_21_315 ();
 FILLCELL_X1 FILLER_0_21_319 ();
 FILLCELL_X4 FILLER_0_21_323 ();
 FILLCELL_X8 FILLER_0_21_330 ();
 FILLCELL_X1 FILLER_0_21_338 ();
 FILLCELL_X2 FILLER_0_21_354 ();
 FILLCELL_X1 FILLER_0_21_362 ();
 FILLCELL_X2 FILLER_0_21_369 ();
 FILLCELL_X1 FILLER_0_21_382 ();
 FILLCELL_X2 FILLER_0_21_394 ();
 FILLCELL_X1 FILLER_0_21_396 ();
 FILLCELL_X1 FILLER_0_21_401 ();
 FILLCELL_X1 FILLER_0_21_417 ();
 FILLCELL_X1 FILLER_0_21_439 ();
 FILLCELL_X4 FILLER_0_22_1 ();
 FILLCELL_X1 FILLER_0_22_5 ();
 FILLCELL_X2 FILLER_0_22_47 ();
 FILLCELL_X2 FILLER_0_22_52 ();
 FILLCELL_X1 FILLER_0_22_54 ();
 FILLCELL_X2 FILLER_0_22_75 ();
 FILLCELL_X2 FILLER_0_22_106 ();
 FILLCELL_X2 FILLER_0_22_124 ();
 FILLCELL_X4 FILLER_0_22_150 ();
 FILLCELL_X1 FILLER_0_22_166 ();
 FILLCELL_X1 FILLER_0_22_169 ();
 FILLCELL_X1 FILLER_0_22_173 ();
 FILLCELL_X2 FILLER_0_22_180 ();
 FILLCELL_X1 FILLER_0_22_185 ();
 FILLCELL_X2 FILLER_0_22_189 ();
 FILLCELL_X1 FILLER_0_22_206 ();
 FILLCELL_X1 FILLER_0_22_217 ();
 FILLCELL_X2 FILLER_0_22_226 ();
 FILLCELL_X2 FILLER_0_22_236 ();
 FILLCELL_X8 FILLER_0_22_241 ();
 FILLCELL_X1 FILLER_0_22_249 ();
 FILLCELL_X8 FILLER_0_22_275 ();
 FILLCELL_X2 FILLER_0_22_283 ();
 FILLCELL_X2 FILLER_0_22_294 ();
 FILLCELL_X4 FILLER_0_22_328 ();
 FILLCELL_X2 FILLER_0_22_332 ();
 FILLCELL_X1 FILLER_0_22_334 ();
 FILLCELL_X1 FILLER_0_22_365 ();
 FILLCELL_X1 FILLER_0_22_382 ();
 FILLCELL_X2 FILLER_0_22_399 ();
 FILLCELL_X2 FILLER_0_22_408 ();
 FILLCELL_X8 FILLER_0_22_419 ();
 FILLCELL_X1 FILLER_0_23_1 ();
 FILLCELL_X1 FILLER_0_23_8 ();
 FILLCELL_X1 FILLER_0_23_13 ();
 FILLCELL_X1 FILLER_0_23_18 ();
 FILLCELL_X1 FILLER_0_23_28 ();
 FILLCELL_X1 FILLER_0_23_33 ();
 FILLCELL_X1 FILLER_0_23_42 ();
 FILLCELL_X1 FILLER_0_23_65 ();
 FILLCELL_X4 FILLER_0_23_83 ();
 FILLCELL_X1 FILLER_0_23_87 ();
 FILLCELL_X1 FILLER_0_23_103 ();
 FILLCELL_X2 FILLER_0_23_123 ();
 FILLCELL_X4 FILLER_0_23_144 ();
 FILLCELL_X1 FILLER_0_23_156 ();
 FILLCELL_X1 FILLER_0_23_177 ();
 FILLCELL_X4 FILLER_0_23_182 ();
 FILLCELL_X2 FILLER_0_23_186 ();
 FILLCELL_X1 FILLER_0_23_188 ();
 FILLCELL_X4 FILLER_0_23_275 ();
 FILLCELL_X2 FILLER_0_23_279 ();
 FILLCELL_X1 FILLER_0_23_281 ();
 FILLCELL_X4 FILLER_0_23_285 ();
 FILLCELL_X8 FILLER_0_23_322 ();
 FILLCELL_X1 FILLER_0_23_336 ();
 FILLCELL_X4 FILLER_0_23_352 ();
 FILLCELL_X2 FILLER_0_23_357 ();
 FILLCELL_X2 FILLER_0_23_408 ();
 FILLCELL_X1 FILLER_0_23_422 ();
 FILLCELL_X8 FILLER_0_23_426 ();
 FILLCELL_X1 FILLER_0_24_25 ();
 FILLCELL_X1 FILLER_0_24_41 ();
 FILLCELL_X2 FILLER_0_24_57 ();
 FILLCELL_X2 FILLER_0_24_65 ();
 FILLCELL_X2 FILLER_0_24_76 ();
 FILLCELL_X1 FILLER_0_24_78 ();
 FILLCELL_X4 FILLER_0_24_85 ();
 FILLCELL_X8 FILLER_0_24_90 ();
 FILLCELL_X2 FILLER_0_24_112 ();
 FILLCELL_X4 FILLER_0_24_122 ();
 FILLCELL_X1 FILLER_0_24_129 ();
 FILLCELL_X2 FILLER_0_24_146 ();
 FILLCELL_X2 FILLER_0_24_175 ();
 FILLCELL_X2 FILLER_0_24_183 ();
 FILLCELL_X1 FILLER_0_24_229 ();
 FILLCELL_X4 FILLER_0_24_233 ();
 FILLCELL_X1 FILLER_0_24_237 ();
 FILLCELL_X4 FILLER_0_24_245 ();
 FILLCELL_X1 FILLER_0_24_249 ();
 FILLCELL_X1 FILLER_0_24_260 ();
 FILLCELL_X2 FILLER_0_24_264 ();
 FILLCELL_X1 FILLER_0_24_266 ();
 FILLCELL_X1 FILLER_0_24_303 ();
 FILLCELL_X1 FILLER_0_24_307 ();
 FILLCELL_X2 FILLER_0_24_311 ();
 FILLCELL_X2 FILLER_0_24_317 ();
 FILLCELL_X1 FILLER_0_24_325 ();
 FILLCELL_X8 FILLER_0_24_349 ();
 FILLCELL_X1 FILLER_0_24_365 ();
 FILLCELL_X2 FILLER_0_24_386 ();
 FILLCELL_X1 FILLER_0_24_391 ();
 FILLCELL_X1 FILLER_0_24_398 ();
 FILLCELL_X1 FILLER_0_24_402 ();
 FILLCELL_X1 FILLER_0_24_407 ();
 FILLCELL_X4 FILLER_0_24_410 ();
 FILLCELL_X1 FILLER_0_24_414 ();
 FILLCELL_X2 FILLER_0_24_438 ();
 FILLCELL_X2 FILLER_0_25_1 ();
 FILLCELL_X1 FILLER_0_25_3 ();
 FILLCELL_X1 FILLER_0_25_27 ();
 FILLCELL_X1 FILLER_0_25_34 ();
 FILLCELL_X1 FILLER_0_25_38 ();
 FILLCELL_X2 FILLER_0_25_46 ();
 FILLCELL_X8 FILLER_0_25_52 ();
 FILLCELL_X4 FILLER_0_25_60 ();
 FILLCELL_X1 FILLER_0_25_64 ();
 FILLCELL_X2 FILLER_0_25_75 ();
 FILLCELL_X8 FILLER_0_25_87 ();
 FILLCELL_X4 FILLER_0_25_95 ();
 FILLCELL_X2 FILLER_0_25_99 ();
 FILLCELL_X1 FILLER_0_25_111 ();
 FILLCELL_X2 FILLER_0_25_122 ();
 FILLCELL_X4 FILLER_0_25_131 ();
 FILLCELL_X1 FILLER_0_25_135 ();
 FILLCELL_X2 FILLER_0_25_164 ();
 FILLCELL_X1 FILLER_0_25_226 ();
 FILLCELL_X4 FILLER_0_25_243 ();
 FILLCELL_X2 FILLER_0_25_247 ();
 FILLCELL_X1 FILLER_0_25_249 ();
 FILLCELL_X1 FILLER_0_25_253 ();
 FILLCELL_X4 FILLER_0_25_258 ();
 FILLCELL_X8 FILLER_0_25_279 ();
 FILLCELL_X2 FILLER_0_25_287 ();
 FILLCELL_X2 FILLER_0_25_296 ();
 FILLCELL_X1 FILLER_0_25_298 ();
 FILLCELL_X2 FILLER_0_25_302 ();
 FILLCELL_X1 FILLER_0_25_304 ();
 FILLCELL_X4 FILLER_0_25_311 ();
 FILLCELL_X1 FILLER_0_25_315 ();
 FILLCELL_X2 FILLER_0_25_318 ();
 FILLCELL_X1 FILLER_0_25_320 ();
 FILLCELL_X2 FILLER_0_25_325 ();
 FILLCELL_X1 FILLER_0_25_327 ();
 FILLCELL_X2 FILLER_0_25_332 ();
 FILLCELL_X1 FILLER_0_25_346 ();
 FILLCELL_X2 FILLER_0_25_357 ();
 FILLCELL_X2 FILLER_0_25_364 ();
 FILLCELL_X2 FILLER_0_25_372 ();
 FILLCELL_X2 FILLER_0_25_380 ();
 FILLCELL_X1 FILLER_0_25_382 ();
 FILLCELL_X1 FILLER_0_25_389 ();
 FILLCELL_X1 FILLER_0_25_396 ();
 FILLCELL_X2 FILLER_0_25_412 ();
 FILLCELL_X1 FILLER_0_25_414 ();
 FILLCELL_X4 FILLER_0_26_1 ();
 FILLCELL_X1 FILLER_0_26_32 ();
 FILLCELL_X2 FILLER_0_26_36 ();
 FILLCELL_X4 FILLER_0_26_44 ();
 FILLCELL_X2 FILLER_0_26_48 ();
 FILLCELL_X2 FILLER_0_26_68 ();
 FILLCELL_X4 FILLER_0_26_111 ();
 FILLCELL_X2 FILLER_0_26_115 ();
 FILLCELL_X1 FILLER_0_26_117 ();
 FILLCELL_X1 FILLER_0_26_130 ();
 FILLCELL_X1 FILLER_0_26_149 ();
 FILLCELL_X2 FILLER_0_26_180 ();
 FILLCELL_X1 FILLER_0_26_200 ();
 FILLCELL_X1 FILLER_0_26_207 ();
 FILLCELL_X2 FILLER_0_26_211 ();
 FILLCELL_X1 FILLER_0_26_213 ();
 FILLCELL_X2 FILLER_0_26_217 ();
 FILLCELL_X4 FILLER_0_26_242 ();
 FILLCELL_X2 FILLER_0_26_246 ();
 FILLCELL_X1 FILLER_0_26_248 ();
 FILLCELL_X1 FILLER_0_26_266 ();
 FILLCELL_X1 FILLER_0_26_268 ();
 FILLCELL_X1 FILLER_0_26_289 ();
 FILLCELL_X1 FILLER_0_26_300 ();
 FILLCELL_X2 FILLER_0_26_305 ();
 FILLCELL_X2 FILLER_0_26_341 ();
 FILLCELL_X2 FILLER_0_26_346 ();
 FILLCELL_X1 FILLER_0_26_348 ();
 FILLCELL_X1 FILLER_0_26_354 ();
 FILLCELL_X2 FILLER_0_26_361 ();
 FILLCELL_X2 FILLER_0_26_371 ();
 FILLCELL_X1 FILLER_0_26_396 ();
 FILLCELL_X1 FILLER_0_26_400 ();
 FILLCELL_X1 FILLER_0_26_409 ();
 FILLCELL_X2 FILLER_0_26_416 ();
 FILLCELL_X1 FILLER_0_26_418 ();
 FILLCELL_X8 FILLER_0_26_425 ();
 FILLCELL_X4 FILLER_0_26_433 ();
 FILLCELL_X2 FILLER_0_26_437 ();
 FILLCELL_X1 FILLER_0_26_439 ();
 FILLCELL_X1 FILLER_0_27_1 ();
 FILLCELL_X4 FILLER_0_27_17 ();
 FILLCELL_X1 FILLER_0_27_25 ();
 FILLCELL_X1 FILLER_0_27_28 ();
 FILLCELL_X2 FILLER_0_27_46 ();
 FILLCELL_X1 FILLER_0_27_48 ();
 FILLCELL_X2 FILLER_0_27_53 ();
 FILLCELL_X4 FILLER_0_27_70 ();
 FILLCELL_X2 FILLER_0_27_80 ();
 FILLCELL_X1 FILLER_0_27_82 ();
 FILLCELL_X8 FILLER_0_27_95 ();
 FILLCELL_X4 FILLER_0_27_103 ();
 FILLCELL_X4 FILLER_0_27_109 ();
 FILLCELL_X1 FILLER_0_27_113 ();
 FILLCELL_X4 FILLER_0_27_124 ();
 FILLCELL_X2 FILLER_0_27_135 ();
 FILLCELL_X1 FILLER_0_27_137 ();
 FILLCELL_X1 FILLER_0_27_145 ();
 FILLCELL_X4 FILLER_0_27_148 ();
 FILLCELL_X1 FILLER_0_27_152 ();
 FILLCELL_X2 FILLER_0_27_170 ();
 FILLCELL_X2 FILLER_0_27_175 ();
 FILLCELL_X1 FILLER_0_27_177 ();
 FILLCELL_X1 FILLER_0_27_179 ();
 FILLCELL_X1 FILLER_0_27_197 ();
 FILLCELL_X1 FILLER_0_27_200 ();
 FILLCELL_X2 FILLER_0_27_205 ();
 FILLCELL_X2 FILLER_0_27_213 ();
 FILLCELL_X2 FILLER_0_27_232 ();
 FILLCELL_X2 FILLER_0_27_237 ();
 FILLCELL_X8 FILLER_0_27_260 ();
 FILLCELL_X1 FILLER_0_27_271 ();
 FILLCELL_X8 FILLER_0_27_275 ();
 FILLCELL_X1 FILLER_0_27_286 ();
 FILLCELL_X4 FILLER_0_27_298 ();
 FILLCELL_X2 FILLER_0_27_302 ();
 FILLCELL_X1 FILLER_0_27_304 ();
 FILLCELL_X2 FILLER_0_27_308 ();
 FILLCELL_X1 FILLER_0_27_310 ();
 FILLCELL_X1 FILLER_0_27_317 ();
 FILLCELL_X1 FILLER_0_27_324 ();
 FILLCELL_X1 FILLER_0_27_328 ();
 FILLCELL_X2 FILLER_0_27_337 ();
 FILLCELL_X2 FILLER_0_27_343 ();
 FILLCELL_X1 FILLER_0_27_345 ();
 FILLCELL_X2 FILLER_0_27_349 ();
 FILLCELL_X1 FILLER_0_27_411 ();
 FILLCELL_X1 FILLER_0_27_417 ();
 FILLCELL_X1 FILLER_0_27_426 ();
 FILLCELL_X8 FILLER_0_27_430 ();
 FILLCELL_X2 FILLER_0_27_438 ();
 FILLCELL_X2 FILLER_0_28_1 ();
 FILLCELL_X1 FILLER_0_28_3 ();
 FILLCELL_X2 FILLER_0_28_16 ();
 FILLCELL_X1 FILLER_0_28_27 ();
 FILLCELL_X1 FILLER_0_28_34 ();
 FILLCELL_X1 FILLER_0_28_42 ();
 FILLCELL_X4 FILLER_0_28_45 ();
 FILLCELL_X1 FILLER_0_28_49 ();
 FILLCELL_X8 FILLER_0_28_53 ();
 FILLCELL_X2 FILLER_0_28_87 ();
 FILLCELL_X4 FILLER_0_28_96 ();
 FILLCELL_X1 FILLER_0_28_100 ();
 FILLCELL_X2 FILLER_0_28_104 ();
 FILLCELL_X1 FILLER_0_28_106 ();
 FILLCELL_X1 FILLER_0_28_124 ();
 FILLCELL_X2 FILLER_0_28_141 ();
 FILLCELL_X1 FILLER_0_28_143 ();
 FILLCELL_X1 FILLER_0_28_150 ();
 FILLCELL_X4 FILLER_0_28_175 ();
 FILLCELL_X2 FILLER_0_28_188 ();
 FILLCELL_X2 FILLER_0_28_208 ();
 FILLCELL_X1 FILLER_0_28_256 ();
 FILLCELL_X4 FILLER_0_28_276 ();
 FILLCELL_X2 FILLER_0_28_280 ();
 FILLCELL_X1 FILLER_0_28_282 ();
 FILLCELL_X4 FILLER_0_28_289 ();
 FILLCELL_X4 FILLER_0_28_300 ();
 FILLCELL_X2 FILLER_0_28_317 ();
 FILLCELL_X8 FILLER_0_28_332 ();
 FILLCELL_X4 FILLER_0_28_379 ();
 FILLCELL_X1 FILLER_0_28_415 ();
 FILLCELL_X4 FILLER_0_28_435 ();
 FILLCELL_X1 FILLER_0_28_439 ();
 FILLCELL_X4 FILLER_0_29_1 ();
 FILLCELL_X2 FILLER_0_29_5 ();
 FILLCELL_X1 FILLER_0_29_7 ();
 FILLCELL_X2 FILLER_0_29_31 ();
 FILLCELL_X4 FILLER_0_29_59 ();
 FILLCELL_X2 FILLER_0_29_63 ();
 FILLCELL_X1 FILLER_0_29_65 ();
 FILLCELL_X4 FILLER_0_29_87 ();
 FILLCELL_X1 FILLER_0_29_91 ();
 FILLCELL_X2 FILLER_0_29_97 ();
 FILLCELL_X1 FILLER_0_29_99 ();
 FILLCELL_X2 FILLER_0_29_106 ();
 FILLCELL_X1 FILLER_0_29_112 ();
 FILLCELL_X1 FILLER_0_29_141 ();
 FILLCELL_X2 FILLER_0_29_172 ();
 FILLCELL_X2 FILLER_0_29_185 ();
 FILLCELL_X8 FILLER_0_29_193 ();
 FILLCELL_X4 FILLER_0_29_201 ();
 FILLCELL_X1 FILLER_0_29_205 ();
 FILLCELL_X1 FILLER_0_29_212 ();
 FILLCELL_X1 FILLER_0_29_216 ();
 FILLCELL_X4 FILLER_0_29_270 ();
 FILLCELL_X1 FILLER_0_29_277 ();
 FILLCELL_X1 FILLER_0_29_288 ();
 FILLCELL_X1 FILLER_0_29_295 ();
 FILLCELL_X1 FILLER_0_29_302 ();
 FILLCELL_X1 FILLER_0_29_306 ();
 FILLCELL_X8 FILLER_0_29_311 ();
 FILLCELL_X1 FILLER_0_29_319 ();
 FILLCELL_X1 FILLER_0_29_350 ();
 FILLCELL_X2 FILLER_0_29_354 ();
 FILLCELL_X1 FILLER_0_29_357 ();
 FILLCELL_X1 FILLER_0_29_364 ();
 FILLCELL_X1 FILLER_0_29_371 ();
 FILLCELL_X1 FILLER_0_29_375 ();
 FILLCELL_X4 FILLER_0_29_379 ();
 FILLCELL_X1 FILLER_0_29_383 ();
 FILLCELL_X2 FILLER_0_29_421 ();
 FILLCELL_X2 FILLER_0_30_1 ();
 FILLCELL_X1 FILLER_0_30_3 ();
 FILLCELL_X2 FILLER_0_30_13 ();
 FILLCELL_X1 FILLER_0_30_15 ();
 FILLCELL_X2 FILLER_0_30_41 ();
 FILLCELL_X2 FILLER_0_30_71 ();
 FILLCELL_X1 FILLER_0_30_93 ();
 FILLCELL_X2 FILLER_0_30_121 ();
 FILLCELL_X1 FILLER_0_30_135 ();
 FILLCELL_X1 FILLER_0_30_142 ();
 FILLCELL_X1 FILLER_0_30_147 ();
 FILLCELL_X2 FILLER_0_30_154 ();
 FILLCELL_X4 FILLER_0_30_162 ();
 FILLCELL_X1 FILLER_0_30_166 ();
 FILLCELL_X1 FILLER_0_30_190 ();
 FILLCELL_X1 FILLER_0_30_197 ();
 FILLCELL_X4 FILLER_0_30_202 ();
 FILLCELL_X1 FILLER_0_30_206 ();
 FILLCELL_X1 FILLER_0_30_217 ();
 FILLCELL_X1 FILLER_0_30_256 ();
 FILLCELL_X1 FILLER_0_30_260 ();
 FILLCELL_X2 FILLER_0_30_298 ();
 FILLCELL_X1 FILLER_0_30_304 ();
 FILLCELL_X4 FILLER_0_30_309 ();
 FILLCELL_X1 FILLER_0_30_313 ();
 FILLCELL_X1 FILLER_0_30_320 ();
 FILLCELL_X2 FILLER_0_30_324 ();
 FILLCELL_X1 FILLER_0_30_326 ();
 FILLCELL_X2 FILLER_0_30_342 ();
 FILLCELL_X8 FILLER_0_30_350 ();
 FILLCELL_X4 FILLER_0_30_358 ();
 FILLCELL_X1 FILLER_0_30_382 ();
 FILLCELL_X1 FILLER_0_30_387 ();
 FILLCELL_X1 FILLER_0_30_391 ();
 FILLCELL_X2 FILLER_0_30_396 ();
 FILLCELL_X1 FILLER_0_30_401 ();
 FILLCELL_X1 FILLER_0_30_406 ();
 FILLCELL_X1 FILLER_0_30_412 ();
 FILLCELL_X2 FILLER_0_30_419 ();
 FILLCELL_X1 FILLER_0_30_435 ();
 FILLCELL_X1 FILLER_0_30_439 ();
 FILLCELL_X8 FILLER_0_31_1 ();
 FILLCELL_X1 FILLER_0_31_13 ();
 FILLCELL_X1 FILLER_0_31_18 ();
 FILLCELL_X1 FILLER_0_31_40 ();
 FILLCELL_X1 FILLER_0_31_47 ();
 FILLCELL_X1 FILLER_0_31_54 ();
 FILLCELL_X2 FILLER_0_31_65 ();
 FILLCELL_X1 FILLER_0_31_67 ();
 FILLCELL_X2 FILLER_0_31_78 ();
 FILLCELL_X1 FILLER_0_31_107 ();
 FILLCELL_X1 FILLER_0_31_123 ();
 FILLCELL_X1 FILLER_0_31_127 ();
 FILLCELL_X2 FILLER_0_31_137 ();
 FILLCELL_X2 FILLER_0_31_149 ();
 FILLCELL_X8 FILLER_0_31_157 ();
 FILLCELL_X4 FILLER_0_31_165 ();
 FILLCELL_X2 FILLER_0_31_169 ();
 FILLCELL_X1 FILLER_0_31_171 ();
 FILLCELL_X1 FILLER_0_31_183 ();
 FILLCELL_X2 FILLER_0_31_193 ();
 FILLCELL_X1 FILLER_0_31_209 ();
 FILLCELL_X1 FILLER_0_31_215 ();
 FILLCELL_X1 FILLER_0_31_219 ();
 FILLCELL_X1 FILLER_0_31_223 ();
 FILLCELL_X2 FILLER_0_31_257 ();
 FILLCELL_X4 FILLER_0_31_271 ();
 FILLCELL_X4 FILLER_0_31_301 ();
 FILLCELL_X2 FILLER_0_31_305 ();
 FILLCELL_X8 FILLER_0_31_324 ();
 FILLCELL_X2 FILLER_0_31_360 ();
 FILLCELL_X1 FILLER_0_31_366 ();
 FILLCELL_X1 FILLER_0_31_372 ();
 FILLCELL_X1 FILLER_0_31_383 ();
 FILLCELL_X1 FILLER_0_31_388 ();
 FILLCELL_X1 FILLER_0_31_395 ();
 FILLCELL_X2 FILLER_0_31_434 ();
 FILLCELL_X1 FILLER_0_31_439 ();
 FILLCELL_X2 FILLER_0_32_1 ();
 FILLCELL_X2 FILLER_0_32_28 ();
 FILLCELL_X1 FILLER_0_32_30 ();
 FILLCELL_X2 FILLER_0_32_35 ();
 FILLCELL_X16 FILLER_0_32_43 ();
 FILLCELL_X8 FILLER_0_32_59 ();
 FILLCELL_X1 FILLER_0_32_67 ();
 FILLCELL_X1 FILLER_0_32_71 ();
 FILLCELL_X2 FILLER_0_32_75 ();
 FILLCELL_X1 FILLER_0_32_77 ();
 FILLCELL_X1 FILLER_0_32_84 ();
 FILLCELL_X8 FILLER_0_32_96 ();
 FILLCELL_X1 FILLER_0_32_108 ();
 FILLCELL_X1 FILLER_0_32_112 ();
 FILLCELL_X1 FILLER_0_32_122 ();
 FILLCELL_X1 FILLER_0_32_132 ();
 FILLCELL_X1 FILLER_0_32_139 ();
 FILLCELL_X1 FILLER_0_32_146 ();
 FILLCELL_X4 FILLER_0_32_163 ();
 FILLCELL_X2 FILLER_0_32_167 ();
 FILLCELL_X1 FILLER_0_32_169 ();
 FILLCELL_X1 FILLER_0_32_173 ();
 FILLCELL_X4 FILLER_0_32_195 ();
 FILLCELL_X2 FILLER_0_32_199 ();
 FILLCELL_X1 FILLER_0_32_201 ();
 FILLCELL_X2 FILLER_0_32_214 ();
 FILLCELL_X1 FILLER_0_32_238 ();
 FILLCELL_X1 FILLER_0_32_243 ();
 FILLCELL_X1 FILLER_0_32_250 ();
 FILLCELL_X1 FILLER_0_32_254 ();
 FILLCELL_X2 FILLER_0_32_259 ();
 FILLCELL_X8 FILLER_0_32_281 ();
 FILLCELL_X1 FILLER_0_32_289 ();
 FILLCELL_X4 FILLER_0_32_299 ();
 FILLCELL_X1 FILLER_0_32_303 ();
 FILLCELL_X16 FILLER_0_32_321 ();
 FILLCELL_X4 FILLER_0_32_339 ();
 FILLCELL_X2 FILLER_0_32_343 ();
 FILLCELL_X4 FILLER_0_32_359 ();
 FILLCELL_X2 FILLER_0_32_363 ();
 FILLCELL_X1 FILLER_0_32_365 ();
 FILLCELL_X1 FILLER_0_32_372 ();
 FILLCELL_X4 FILLER_0_32_388 ();
 FILLCELL_X2 FILLER_0_32_392 ();
 FILLCELL_X2 FILLER_0_32_397 ();
 FILLCELL_X1 FILLER_0_32_402 ();
 FILLCELL_X1 FILLER_0_32_409 ();
 FILLCELL_X1 FILLER_0_32_414 ();
 FILLCELL_X1 FILLER_0_32_425 ();
 FILLCELL_X1 FILLER_0_32_432 ();
 FILLCELL_X1 FILLER_0_33_12 ();
 FILLCELL_X2 FILLER_0_33_25 ();
 FILLCELL_X1 FILLER_0_33_27 ();
 FILLCELL_X2 FILLER_0_33_47 ();
 FILLCELL_X1 FILLER_0_33_66 ();
 FILLCELL_X1 FILLER_0_33_94 ();
 FILLCELL_X1 FILLER_0_33_101 ();
 FILLCELL_X8 FILLER_0_33_119 ();
 FILLCELL_X1 FILLER_0_33_139 ();
 FILLCELL_X1 FILLER_0_33_147 ();
 FILLCELL_X4 FILLER_0_33_154 ();
 FILLCELL_X4 FILLER_0_33_196 ();
 FILLCELL_X2 FILLER_0_33_226 ();
 FILLCELL_X1 FILLER_0_33_232 ();
 FILLCELL_X1 FILLER_0_33_243 ();
 FILLCELL_X1 FILLER_0_33_247 ();
 FILLCELL_X2 FILLER_0_33_257 ();
 FILLCELL_X1 FILLER_0_33_287 ();
 FILLCELL_X2 FILLER_0_33_292 ();
 FILLCELL_X2 FILLER_0_33_300 ();
 FILLCELL_X2 FILLER_0_33_308 ();
 FILLCELL_X1 FILLER_0_33_310 ();
 FILLCELL_X4 FILLER_0_33_315 ();
 FILLCELL_X2 FILLER_0_33_319 ();
 FILLCELL_X1 FILLER_0_33_321 ();
 FILLCELL_X1 FILLER_0_33_328 ();
 FILLCELL_X8 FILLER_0_33_337 ();
 FILLCELL_X4 FILLER_0_33_345 ();
 FILLCELL_X2 FILLER_0_33_354 ();
 FILLCELL_X2 FILLER_0_33_387 ();
 FILLCELL_X1 FILLER_0_33_389 ();
 FILLCELL_X4 FILLER_0_33_397 ();
 FILLCELL_X2 FILLER_0_33_401 ();
 FILLCELL_X1 FILLER_0_33_403 ();
 FILLCELL_X1 FILLER_0_33_407 ();
 FILLCELL_X1 FILLER_0_33_414 ();
 FILLCELL_X4 FILLER_0_33_430 ();
 FILLCELL_X2 FILLER_0_33_437 ();
 FILLCELL_X1 FILLER_0_33_439 ();
 FILLCELL_X1 FILLER_0_34_16 ();
 FILLCELL_X1 FILLER_0_34_21 ();
 FILLCELL_X1 FILLER_0_34_34 ();
 FILLCELL_X1 FILLER_0_34_41 ();
 FILLCELL_X1 FILLER_0_34_45 ();
 FILLCELL_X4 FILLER_0_34_60 ();
 FILLCELL_X1 FILLER_0_34_64 ();
 FILLCELL_X4 FILLER_0_34_77 ();
 FILLCELL_X2 FILLER_0_34_81 ();
 FILLCELL_X2 FILLER_0_34_87 ();
 FILLCELL_X8 FILLER_0_34_93 ();
 FILLCELL_X4 FILLER_0_34_101 ();
 FILLCELL_X1 FILLER_0_34_105 ();
 FILLCELL_X2 FILLER_0_34_117 ();
 FILLCELL_X1 FILLER_0_34_161 ();
 FILLCELL_X4 FILLER_0_34_168 ();
 FILLCELL_X2 FILLER_0_34_172 ();
 FILLCELL_X1 FILLER_0_34_174 ();
 FILLCELL_X2 FILLER_0_34_179 ();
 FILLCELL_X1 FILLER_0_34_188 ();
 FILLCELL_X2 FILLER_0_34_212 ();
 FILLCELL_X1 FILLER_0_34_214 ();
 FILLCELL_X2 FILLER_0_34_233 ();
 FILLCELL_X1 FILLER_0_34_235 ();
 FILLCELL_X1 FILLER_0_34_254 ();
 FILLCELL_X2 FILLER_0_34_265 ();
 FILLCELL_X2 FILLER_0_34_268 ();
 FILLCELL_X1 FILLER_0_34_285 ();
 FILLCELL_X1 FILLER_0_34_289 ();
 FILLCELL_X1 FILLER_0_34_296 ();
 FILLCELL_X1 FILLER_0_34_300 ();
 FILLCELL_X1 FILLER_0_34_318 ();
 FILLCELL_X1 FILLER_0_34_322 ();
 FILLCELL_X2 FILLER_0_34_327 ();
 FILLCELL_X2 FILLER_0_34_348 ();
 FILLCELL_X2 FILLER_0_34_381 ();
 FILLCELL_X1 FILLER_0_34_400 ();
 FILLCELL_X2 FILLER_0_34_427 ();
 FILLCELL_X8 FILLER_0_34_432 ();
 FILLCELL_X1 FILLER_0_35_1 ();
 FILLCELL_X2 FILLER_0_35_12 ();
 FILLCELL_X2 FILLER_0_35_19 ();
 FILLCELL_X1 FILLER_0_35_21 ();
 FILLCELL_X2 FILLER_0_35_34 ();
 FILLCELL_X1 FILLER_0_35_42 ();
 FILLCELL_X1 FILLER_0_35_53 ();
 FILLCELL_X4 FILLER_0_35_61 ();
 FILLCELL_X2 FILLER_0_35_65 ();
 FILLCELL_X1 FILLER_0_35_70 ();
 FILLCELL_X2 FILLER_0_35_86 ();
 FILLCELL_X1 FILLER_0_35_95 ();
 FILLCELL_X1 FILLER_0_35_102 ();
 FILLCELL_X1 FILLER_0_35_106 ();
 FILLCELL_X1 FILLER_0_35_113 ();
 FILLCELL_X2 FILLER_0_35_141 ();
 FILLCELL_X2 FILLER_0_35_167 ();
 FILLCELL_X1 FILLER_0_35_179 ();
 FILLCELL_X1 FILLER_0_35_193 ();
 FILLCELL_X4 FILLER_0_35_197 ();
 FILLCELL_X1 FILLER_0_35_201 ();
 FILLCELL_X2 FILLER_0_35_205 ();
 FILLCELL_X2 FILLER_0_35_220 ();
 FILLCELL_X1 FILLER_0_35_222 ();
 FILLCELL_X1 FILLER_0_35_229 ();
 FILLCELL_X2 FILLER_0_35_259 ();
 FILLCELL_X1 FILLER_0_35_264 ();
 FILLCELL_X1 FILLER_0_35_271 ();
 FILLCELL_X4 FILLER_0_35_288 ();
 FILLCELL_X8 FILLER_0_35_299 ();
 FILLCELL_X4 FILLER_0_35_310 ();
 FILLCELL_X1 FILLER_0_35_331 ();
 FILLCELL_X2 FILLER_0_35_337 ();
 FILLCELL_X2 FILLER_0_35_346 ();
 FILLCELL_X2 FILLER_0_35_357 ();
 FILLCELL_X1 FILLER_0_35_359 ();
 FILLCELL_X4 FILLER_0_35_370 ();
 FILLCELL_X2 FILLER_0_35_374 ();
 FILLCELL_X2 FILLER_0_35_379 ();
 FILLCELL_X1 FILLER_0_35_381 ();
 FILLCELL_X1 FILLER_0_35_403 ();
 FILLCELL_X2 FILLER_0_35_427 ();
 FILLCELL_X1 FILLER_0_35_429 ();
 FILLCELL_X2 FILLER_0_36_1 ();
 FILLCELL_X8 FILLER_0_36_15 ();
 FILLCELL_X4 FILLER_0_36_23 ();
 FILLCELL_X4 FILLER_0_36_33 ();
 FILLCELL_X2 FILLER_0_36_37 ();
 FILLCELL_X2 FILLER_0_36_55 ();
 FILLCELL_X4 FILLER_0_36_61 ();
 FILLCELL_X1 FILLER_0_36_131 ();
 FILLCELL_X1 FILLER_0_36_136 ();
 FILLCELL_X1 FILLER_0_36_146 ();
 FILLCELL_X1 FILLER_0_36_150 ();
 FILLCELL_X1 FILLER_0_36_154 ();
 FILLCELL_X1 FILLER_0_36_159 ();
 FILLCELL_X1 FILLER_0_36_175 ();
 FILLCELL_X1 FILLER_0_36_179 ();
 FILLCELL_X2 FILLER_0_36_190 ();
 FILLCELL_X2 FILLER_0_36_209 ();
 FILLCELL_X4 FILLER_0_36_228 ();
 FILLCELL_X1 FILLER_0_36_241 ();
 FILLCELL_X1 FILLER_0_36_245 ();
 FILLCELL_X1 FILLER_0_36_255 ();
 FILLCELL_X2 FILLER_0_36_262 ();
 FILLCELL_X2 FILLER_0_36_299 ();
 FILLCELL_X8 FILLER_0_36_313 ();
 FILLCELL_X16 FILLER_0_36_331 ();
 FILLCELL_X2 FILLER_0_36_369 ();
 FILLCELL_X2 FILLER_0_36_380 ();
 FILLCELL_X1 FILLER_0_36_382 ();
 FILLCELL_X2 FILLER_0_36_417 ();
 FILLCELL_X1 FILLER_0_36_422 ();
 FILLCELL_X2 FILLER_0_37_16 ();
 FILLCELL_X1 FILLER_0_37_22 ();
 FILLCELL_X2 FILLER_0_37_29 ();
 FILLCELL_X8 FILLER_0_37_41 ();
 FILLCELL_X4 FILLER_0_37_49 ();
 FILLCELL_X2 FILLER_0_37_78 ();
 FILLCELL_X1 FILLER_0_37_106 ();
 FILLCELL_X2 FILLER_0_37_111 ();
 FILLCELL_X4 FILLER_0_37_140 ();
 FILLCELL_X2 FILLER_0_37_144 ();
 FILLCELL_X2 FILLER_0_37_176 ();
 FILLCELL_X1 FILLER_0_37_179 ();
 FILLCELL_X1 FILLER_0_37_187 ();
 FILLCELL_X1 FILLER_0_37_191 ();
 FILLCELL_X2 FILLER_0_37_211 ();
 FILLCELL_X1 FILLER_0_37_219 ();
 FILLCELL_X1 FILLER_0_37_223 ();
 FILLCELL_X1 FILLER_0_37_241 ();
 FILLCELL_X2 FILLER_0_37_248 ();
 FILLCELL_X2 FILLER_0_37_263 ();
 FILLCELL_X1 FILLER_0_37_265 ();
 FILLCELL_X4 FILLER_0_37_293 ();
 FILLCELL_X2 FILLER_0_37_300 ();
 FILLCELL_X1 FILLER_0_37_315 ();
 FILLCELL_X4 FILLER_0_37_319 ();
 FILLCELL_X1 FILLER_0_37_323 ();
 FILLCELL_X1 FILLER_0_37_341 ();
 FILLCELL_X1 FILLER_0_37_348 ();
 FILLCELL_X4 FILLER_0_37_352 ();
 FILLCELL_X4 FILLER_0_37_357 ();
 FILLCELL_X1 FILLER_0_37_395 ();
 FILLCELL_X1 FILLER_0_37_405 ();
 FILLCELL_X2 FILLER_0_37_424 ();
 FILLCELL_X4 FILLER_0_37_429 ();
 FILLCELL_X1 FILLER_0_37_433 ();
 FILLCELL_X4 FILLER_0_38_1 ();
 FILLCELL_X1 FILLER_0_38_12 ();
 FILLCELL_X1 FILLER_0_38_30 ();
 FILLCELL_X1 FILLER_0_38_35 ();
 FILLCELL_X1 FILLER_0_38_39 ();
 FILLCELL_X1 FILLER_0_38_43 ();
 FILLCELL_X2 FILLER_0_38_48 ();
 FILLCELL_X1 FILLER_0_38_53 ();
 FILLCELL_X1 FILLER_0_38_108 ();
 FILLCELL_X4 FILLER_0_38_130 ();
 FILLCELL_X2 FILLER_0_38_134 ();
 FILLCELL_X2 FILLER_0_38_140 ();
 FILLCELL_X1 FILLER_0_38_201 ();
 FILLCELL_X1 FILLER_0_38_205 ();
 FILLCELL_X1 FILLER_0_38_216 ();
 FILLCELL_X2 FILLER_0_38_220 ();
 FILLCELL_X2 FILLER_0_38_228 ();
 FILLCELL_X1 FILLER_0_38_230 ();
 FILLCELL_X2 FILLER_0_38_257 ();
 FILLCELL_X2 FILLER_0_38_265 ();
 FILLCELL_X1 FILLER_0_38_300 ();
 FILLCELL_X1 FILLER_0_38_358 ();
 FILLCELL_X1 FILLER_0_38_364 ();
 FILLCELL_X1 FILLER_0_38_373 ();
 FILLCELL_X1 FILLER_0_38_380 ();
 FILLCELL_X1 FILLER_0_38_387 ();
 FILLCELL_X1 FILLER_0_38_396 ();
 FILLCELL_X1 FILLER_0_38_424 ();
 FILLCELL_X2 FILLER_0_38_434 ();
 FILLCELL_X1 FILLER_0_38_439 ();
 FILLCELL_X1 FILLER_0_39_37 ();
 FILLCELL_X1 FILLER_0_39_41 ();
 FILLCELL_X4 FILLER_0_39_48 ();
 FILLCELL_X1 FILLER_0_39_52 ();
 FILLCELL_X2 FILLER_0_39_59 ();
 FILLCELL_X1 FILLER_0_39_65 ();
 FILLCELL_X4 FILLER_0_39_72 ();
 FILLCELL_X1 FILLER_0_39_80 ();
 FILLCELL_X2 FILLER_0_39_91 ();
 FILLCELL_X2 FILLER_0_39_102 ();
 FILLCELL_X1 FILLER_0_39_104 ();
 FILLCELL_X4 FILLER_0_39_108 ();
 FILLCELL_X1 FILLER_0_39_112 ();
 FILLCELL_X1 FILLER_0_39_116 ();
 FILLCELL_X2 FILLER_0_39_123 ();
 FILLCELL_X1 FILLER_0_39_201 ();
 FILLCELL_X4 FILLER_0_39_226 ();
 FILLCELL_X8 FILLER_0_39_250 ();
 FILLCELL_X2 FILLER_0_39_264 ();
 FILLCELL_X1 FILLER_0_39_266 ();
 FILLCELL_X4 FILLER_0_39_304 ();
 FILLCELL_X1 FILLER_0_39_324 ();
 FILLCELL_X8 FILLER_0_39_328 ();
 FILLCELL_X4 FILLER_0_39_336 ();
 FILLCELL_X2 FILLER_0_39_343 ();
 FILLCELL_X1 FILLER_0_39_345 ();
 FILLCELL_X1 FILLER_0_39_355 ();
 FILLCELL_X2 FILLER_0_39_374 ();
 FILLCELL_X1 FILLER_0_39_376 ();
 FILLCELL_X1 FILLER_0_39_428 ();
 FILLCELL_X1 FILLER_0_39_435 ();
 FILLCELL_X4 FILLER_0_40_1 ();
 FILLCELL_X1 FILLER_0_40_5 ();
 FILLCELL_X1 FILLER_0_40_17 ();
 FILLCELL_X1 FILLER_0_40_20 ();
 FILLCELL_X1 FILLER_0_40_24 ();
 FILLCELL_X2 FILLER_0_40_28 ();
 FILLCELL_X1 FILLER_0_40_53 ();
 FILLCELL_X2 FILLER_0_40_57 ();
 FILLCELL_X1 FILLER_0_40_59 ();
 FILLCELL_X2 FILLER_0_40_63 ();
 FILLCELL_X2 FILLER_0_40_99 ();
 FILLCELL_X1 FILLER_0_40_104 ();
 FILLCELL_X2 FILLER_0_40_121 ();
 FILLCELL_X1 FILLER_0_40_155 ();
 FILLCELL_X1 FILLER_0_40_165 ();
 FILLCELL_X1 FILLER_0_40_206 ();
 FILLCELL_X1 FILLER_0_40_213 ();
 FILLCELL_X1 FILLER_0_40_224 ();
 FILLCELL_X1 FILLER_0_40_234 ();
 FILLCELL_X4 FILLER_0_40_238 ();
 FILLCELL_X1 FILLER_0_40_242 ();
 FILLCELL_X4 FILLER_0_40_250 ();
 FILLCELL_X1 FILLER_0_40_254 ();
 FILLCELL_X2 FILLER_0_40_286 ();
 FILLCELL_X1 FILLER_0_40_301 ();
 FILLCELL_X2 FILLER_0_40_334 ();
 FILLCELL_X4 FILLER_0_40_360 ();
 FILLCELL_X2 FILLER_0_40_364 ();
 FILLCELL_X1 FILLER_0_40_366 ();
 FILLCELL_X1 FILLER_0_40_369 ();
 FILLCELL_X2 FILLER_0_40_373 ();
 FILLCELL_X1 FILLER_0_40_378 ();
 FILLCELL_X1 FILLER_0_40_382 ();
 FILLCELL_X1 FILLER_0_40_389 ();
 FILLCELL_X1 FILLER_0_40_394 ();
 FILLCELL_X1 FILLER_0_40_399 ();
 FILLCELL_X1 FILLER_0_40_410 ();
 FILLCELL_X2 FILLER_0_40_427 ();
 FILLCELL_X4 FILLER_0_40_433 ();
 FILLCELL_X4 FILLER_0_41_1 ();
 FILLCELL_X2 FILLER_0_41_5 ();
 FILLCELL_X1 FILLER_0_41_25 ();
 FILLCELL_X4 FILLER_0_41_41 ();
 FILLCELL_X1 FILLER_0_41_51 ();
 FILLCELL_X2 FILLER_0_41_58 ();
 FILLCELL_X2 FILLER_0_41_82 ();
 FILLCELL_X1 FILLER_0_41_109 ();
 FILLCELL_X2 FILLER_0_41_113 ();
 FILLCELL_X1 FILLER_0_41_115 ();
 FILLCELL_X2 FILLER_0_41_149 ();
 FILLCELL_X2 FILLER_0_41_167 ();
 FILLCELL_X1 FILLER_0_41_204 ();
 FILLCELL_X1 FILLER_0_41_214 ();
 FILLCELL_X1 FILLER_0_41_218 ();
 FILLCELL_X4 FILLER_0_41_229 ();
 FILLCELL_X1 FILLER_0_41_233 ();
 FILLCELL_X4 FILLER_0_41_238 ();
 FILLCELL_X2 FILLER_0_41_242 ();
 FILLCELL_X1 FILLER_0_41_250 ();
 FILLCELL_X1 FILLER_0_41_274 ();
 FILLCELL_X1 FILLER_0_41_278 ();
 FILLCELL_X1 FILLER_0_41_292 ();
 FILLCELL_X1 FILLER_0_41_299 ();
 FILLCELL_X1 FILLER_0_41_306 ();
 FILLCELL_X8 FILLER_0_41_326 ();
 FILLCELL_X4 FILLER_0_41_334 ();
 FILLCELL_X1 FILLER_0_41_338 ();
 FILLCELL_X1 FILLER_0_41_363 ();
 FILLCELL_X1 FILLER_0_41_370 ();
 FILLCELL_X1 FILLER_0_41_377 ();
 FILLCELL_X1 FILLER_0_41_384 ();
 FILLCELL_X2 FILLER_0_41_389 ();
 FILLCELL_X2 FILLER_0_41_395 ();
 FILLCELL_X1 FILLER_0_41_403 ();
 FILLCELL_X2 FILLER_0_41_408 ();
 FILLCELL_X1 FILLER_0_41_410 ();
 FILLCELL_X2 FILLER_0_41_421 ();
 FILLCELL_X1 FILLER_0_41_439 ();
 FILLCELL_X1 FILLER_0_42_1 ();
 FILLCELL_X2 FILLER_0_42_17 ();
 FILLCELL_X1 FILLER_0_42_19 ();
 FILLCELL_X1 FILLER_0_42_26 ();
 FILLCELL_X1 FILLER_0_42_34 ();
 FILLCELL_X1 FILLER_0_42_39 ();
 FILLCELL_X1 FILLER_0_42_43 ();
 FILLCELL_X1 FILLER_0_42_47 ();
 FILLCELL_X1 FILLER_0_42_51 ();
 FILLCELL_X1 FILLER_0_42_58 ();
 FILLCELL_X2 FILLER_0_42_76 ();
 FILLCELL_X1 FILLER_0_42_84 ();
 FILLCELL_X2 FILLER_0_42_109 ();
 FILLCELL_X1 FILLER_0_42_131 ();
 FILLCELL_X1 FILLER_0_42_135 ();
 FILLCELL_X1 FILLER_0_42_153 ();
 FILLCELL_X1 FILLER_0_42_171 ();
 FILLCELL_X1 FILLER_0_42_178 ();
 FILLCELL_X1 FILLER_0_42_182 ();
 FILLCELL_X1 FILLER_0_42_186 ();
 FILLCELL_X1 FILLER_0_42_205 ();
 FILLCELL_X1 FILLER_0_42_209 ();
 FILLCELL_X2 FILLER_0_42_231 ();
 FILLCELL_X4 FILLER_0_42_256 ();
 FILLCELL_X2 FILLER_0_42_260 ();
 FILLCELL_X1 FILLER_0_42_266 ();
 FILLCELL_X1 FILLER_0_42_274 ();
 FILLCELL_X1 FILLER_0_42_281 ();
 FILLCELL_X1 FILLER_0_42_308 ();
 FILLCELL_X1 FILLER_0_42_325 ();
 FILLCELL_X2 FILLER_0_42_338 ();
 FILLCELL_X1 FILLER_0_42_347 ();
 FILLCELL_X1 FILLER_0_42_406 ();
 FILLCELL_X1 FILLER_0_42_410 ();
 FILLCELL_X1 FILLER_0_42_419 ();
 FILLCELL_X2 FILLER_0_42_424 ();
 FILLCELL_X1 FILLER_0_42_430 ();
 FILLCELL_X1 FILLER_0_42_434 ();
 FILLCELL_X4 FILLER_0_43_1 ();
 FILLCELL_X1 FILLER_0_43_21 ();
 FILLCELL_X1 FILLER_0_43_28 ();
 FILLCELL_X4 FILLER_0_43_35 ();
 FILLCELL_X1 FILLER_0_43_48 ();
 FILLCELL_X1 FILLER_0_43_52 ();
 FILLCELL_X1 FILLER_0_43_60 ();
 FILLCELL_X4 FILLER_0_43_64 ();
 FILLCELL_X2 FILLER_0_43_68 ();
 FILLCELL_X1 FILLER_0_43_70 ();
 FILLCELL_X2 FILLER_0_43_85 ();
 FILLCELL_X2 FILLER_0_43_107 ();
 FILLCELL_X1 FILLER_0_43_115 ();
 FILLCELL_X1 FILLER_0_43_125 ();
 FILLCELL_X1 FILLER_0_43_174 ();
 FILLCELL_X1 FILLER_0_43_185 ();
 FILLCELL_X2 FILLER_0_43_191 ();
 FILLCELL_X2 FILLER_0_43_220 ();
 FILLCELL_X8 FILLER_0_43_238 ();
 FILLCELL_X4 FILLER_0_43_246 ();
 FILLCELL_X2 FILLER_0_43_287 ();
 FILLCELL_X2 FILLER_0_43_308 ();
 FILLCELL_X2 FILLER_0_43_326 ();
 FILLCELL_X1 FILLER_0_43_338 ();
 FILLCELL_X1 FILLER_0_43_348 ();
 FILLCELL_X1 FILLER_0_43_380 ();
 FILLCELL_X2 FILLER_0_43_387 ();
 FILLCELL_X2 FILLER_0_43_395 ();
 FILLCELL_X1 FILLER_0_43_397 ();
 FILLCELL_X1 FILLER_0_43_401 ();
 FILLCELL_X1 FILLER_0_43_408 ();
 FILLCELL_X1 FILLER_0_43_413 ();
 FILLCELL_X1 FILLER_0_43_417 ();
 FILLCELL_X4 FILLER_0_44_1 ();
 FILLCELL_X2 FILLER_0_44_5 ();
 FILLCELL_X1 FILLER_0_44_24 ();
 FILLCELL_X1 FILLER_0_44_28 ();
 FILLCELL_X1 FILLER_0_44_32 ();
 FILLCELL_X4 FILLER_0_44_62 ();
 FILLCELL_X2 FILLER_0_44_66 ();
 FILLCELL_X2 FILLER_0_44_74 ();
 FILLCELL_X1 FILLER_0_44_79 ();
 FILLCELL_X1 FILLER_0_44_107 ();
 FILLCELL_X2 FILLER_0_44_111 ();
 FILLCELL_X8 FILLER_0_44_119 ();
 FILLCELL_X1 FILLER_0_44_127 ();
 FILLCELL_X1 FILLER_0_44_170 ();
 FILLCELL_X2 FILLER_0_44_186 ();
 FILLCELL_X1 FILLER_0_44_197 ();
 FILLCELL_X1 FILLER_0_44_201 ();
 FILLCELL_X1 FILLER_0_44_206 ();
 FILLCELL_X1 FILLER_0_44_210 ();
 FILLCELL_X1 FILLER_0_44_214 ();
 FILLCELL_X4 FILLER_0_44_221 ();
 FILLCELL_X1 FILLER_0_44_225 ();
 FILLCELL_X2 FILLER_0_44_247 ();
 FILLCELL_X2 FILLER_0_44_252 ();
 FILLCELL_X1 FILLER_0_44_254 ();
 FILLCELL_X2 FILLER_0_44_278 ();
 FILLCELL_X2 FILLER_0_44_301 ();
 FILLCELL_X1 FILLER_0_44_303 ();
 FILLCELL_X2 FILLER_0_44_310 ();
 FILLCELL_X2 FILLER_0_44_318 ();
 FILLCELL_X1 FILLER_0_44_341 ();
 FILLCELL_X2 FILLER_0_44_346 ();
 FILLCELL_X1 FILLER_0_44_348 ();
 FILLCELL_X1 FILLER_0_44_361 ();
 FILLCELL_X2 FILLER_0_44_365 ();
 FILLCELL_X2 FILLER_0_44_373 ();
 FILLCELL_X1 FILLER_0_44_375 ();
 FILLCELL_X4 FILLER_0_44_386 ();
 FILLCELL_X4 FILLER_0_44_404 ();
 FILLCELL_X2 FILLER_0_44_408 ();
 FILLCELL_X1 FILLER_0_44_410 ();
 FILLCELL_X1 FILLER_0_44_420 ();
 FILLCELL_X1 FILLER_0_44_427 ();
 FILLCELL_X1 FILLER_0_44_431 ();
 FILLCELL_X4 FILLER_0_44_435 ();
 FILLCELL_X1 FILLER_0_44_439 ();
 FILLCELL_X8 FILLER_0_45_1 ();
 FILLCELL_X2 FILLER_0_45_16 ();
 FILLCELL_X1 FILLER_0_45_18 ();
 FILLCELL_X2 FILLER_0_45_23 ();
 FILLCELL_X2 FILLER_0_45_40 ();
 FILLCELL_X1 FILLER_0_45_51 ();
 FILLCELL_X2 FILLER_0_45_64 ();
 FILLCELL_X2 FILLER_0_45_69 ();
 FILLCELL_X1 FILLER_0_45_94 ();
 FILLCELL_X4 FILLER_0_45_105 ();
 FILLCELL_X2 FILLER_0_45_122 ();
 FILLCELL_X1 FILLER_0_45_127 ();
 FILLCELL_X1 FILLER_0_45_141 ();
 FILLCELL_X1 FILLER_0_45_179 ();
 FILLCELL_X1 FILLER_0_45_186 ();
 FILLCELL_X1 FILLER_0_45_194 ();
 FILLCELL_X1 FILLER_0_45_208 ();
 FILLCELL_X1 FILLER_0_45_215 ();
 FILLCELL_X4 FILLER_0_45_220 ();
 FILLCELL_X1 FILLER_0_45_224 ();
 FILLCELL_X2 FILLER_0_45_250 ();
 FILLCELL_X1 FILLER_0_45_298 ();
 FILLCELL_X1 FILLER_0_45_306 ();
 FILLCELL_X8 FILLER_0_45_360 ();
 FILLCELL_X4 FILLER_0_45_368 ();
 FILLCELL_X2 FILLER_0_45_421 ();
 FILLCELL_X2 FILLER_0_45_435 ();
 FILLCELL_X2 FILLER_0_46_1 ();
 FILLCELL_X1 FILLER_0_46_3 ();
 FILLCELL_X4 FILLER_0_46_49 ();
 FILLCELL_X2 FILLER_0_46_53 ();
 FILLCELL_X2 FILLER_0_46_64 ();
 FILLCELL_X1 FILLER_0_46_66 ();
 FILLCELL_X4 FILLER_0_46_73 ();
 FILLCELL_X1 FILLER_0_46_77 ();
 FILLCELL_X2 FILLER_0_46_80 ();
 FILLCELL_X1 FILLER_0_46_82 ();
 FILLCELL_X4 FILLER_0_46_120 ();
 FILLCELL_X1 FILLER_0_46_127 ();
 FILLCELL_X1 FILLER_0_46_148 ();
 FILLCELL_X1 FILLER_0_46_184 ();
 FILLCELL_X2 FILLER_0_46_210 ();
 FILLCELL_X1 FILLER_0_46_215 ();
 FILLCELL_X1 FILLER_0_46_222 ();
 FILLCELL_X4 FILLER_0_46_260 ();
 FILLCELL_X2 FILLER_0_46_264 ();
 FILLCELL_X1 FILLER_0_46_266 ();
 FILLCELL_X1 FILLER_0_46_310 ();
 FILLCELL_X2 FILLER_0_46_326 ();
 FILLCELL_X1 FILLER_0_46_328 ();
 FILLCELL_X1 FILLER_0_46_333 ();
 FILLCELL_X2 FILLER_0_46_337 ();
 FILLCELL_X2 FILLER_0_46_348 ();
 FILLCELL_X1 FILLER_0_46_356 ();
 FILLCELL_X1 FILLER_0_46_363 ();
 FILLCELL_X1 FILLER_0_46_370 ();
 FILLCELL_X1 FILLER_0_46_374 ();
 FILLCELL_X1 FILLER_0_46_377 ();
 FILLCELL_X1 FILLER_0_46_383 ();
 FILLCELL_X1 FILLER_0_46_388 ();
 FILLCELL_X1 FILLER_0_46_393 ();
 FILLCELL_X4 FILLER_0_46_399 ();
 FILLCELL_X2 FILLER_0_46_403 ();
 FILLCELL_X1 FILLER_0_46_433 ();
 FILLCELL_X4 FILLER_0_47_1 ();
 FILLCELL_X2 FILLER_0_47_5 ();
 FILLCELL_X4 FILLER_0_47_51 ();
 FILLCELL_X2 FILLER_0_47_55 ();
 FILLCELL_X2 FILLER_0_47_63 ();
 FILLCELL_X1 FILLER_0_47_65 ();
 FILLCELL_X2 FILLER_0_47_72 ();
 FILLCELL_X1 FILLER_0_47_74 ();
 FILLCELL_X2 FILLER_0_47_78 ();
 FILLCELL_X1 FILLER_0_47_90 ();
 FILLCELL_X1 FILLER_0_47_102 ();
 FILLCELL_X1 FILLER_0_47_137 ();
 FILLCELL_X2 FILLER_0_47_201 ();
 FILLCELL_X1 FILLER_0_47_203 ();
 FILLCELL_X2 FILLER_0_47_213 ();
 FILLCELL_X1 FILLER_0_47_221 ();
 FILLCELL_X1 FILLER_0_47_228 ();
 FILLCELL_X1 FILLER_0_47_243 ();
 FILLCELL_X1 FILLER_0_47_256 ();
 FILLCELL_X8 FILLER_0_47_260 ();
 FILLCELL_X4 FILLER_0_47_268 ();
 FILLCELL_X2 FILLER_0_47_272 ();
 FILLCELL_X1 FILLER_0_47_280 ();
 FILLCELL_X1 FILLER_0_47_284 ();
 FILLCELL_X1 FILLER_0_47_291 ();
 FILLCELL_X1 FILLER_0_47_296 ();
 FILLCELL_X1 FILLER_0_47_309 ();
 FILLCELL_X2 FILLER_0_47_342 ();
 FILLCELL_X1 FILLER_0_47_344 ();
 FILLCELL_X1 FILLER_0_47_357 ();
 FILLCELL_X1 FILLER_0_47_364 ();
 FILLCELL_X2 FILLER_0_47_369 ();
 FILLCELL_X1 FILLER_0_47_376 ();
 FILLCELL_X1 FILLER_0_47_379 ();
 FILLCELL_X1 FILLER_0_47_387 ();
 FILLCELL_X2 FILLER_0_47_402 ();
 FILLCELL_X4 FILLER_0_47_436 ();
 FILLCELL_X1 FILLER_0_48_4 ();
 FILLCELL_X4 FILLER_0_48_8 ();
 FILLCELL_X1 FILLER_0_48_26 ();
 FILLCELL_X2 FILLER_0_48_35 ();
 FILLCELL_X4 FILLER_0_48_43 ();
 FILLCELL_X2 FILLER_0_48_47 ();
 FILLCELL_X1 FILLER_0_48_49 ();
 FILLCELL_X4 FILLER_0_48_53 ();
 FILLCELL_X2 FILLER_0_48_73 ();
 FILLCELL_X8 FILLER_0_48_81 ();
 FILLCELL_X2 FILLER_0_48_105 ();
 FILLCELL_X2 FILLER_0_48_110 ();
 FILLCELL_X1 FILLER_0_48_138 ();
 FILLCELL_X1 FILLER_0_48_164 ();
 FILLCELL_X2 FILLER_0_48_168 ();
 FILLCELL_X1 FILLER_0_48_170 ();
 FILLCELL_X2 FILLER_0_48_196 ();
 FILLCELL_X1 FILLER_0_48_204 ();
 FILLCELL_X1 FILLER_0_48_215 ();
 FILLCELL_X1 FILLER_0_48_234 ();
 FILLCELL_X2 FILLER_0_48_239 ();
 FILLCELL_X2 FILLER_0_48_245 ();
 FILLCELL_X2 FILLER_0_48_268 ();
 FILLCELL_X8 FILLER_0_48_276 ();
 FILLCELL_X1 FILLER_0_48_310 ();
 FILLCELL_X1 FILLER_0_48_315 ();
 FILLCELL_X1 FILLER_0_48_322 ();
 FILLCELL_X1 FILLER_0_48_332 ();
 FILLCELL_X2 FILLER_0_48_337 ();
 FILLCELL_X2 FILLER_0_48_356 ();
 FILLCELL_X2 FILLER_0_48_361 ();
 FILLCELL_X2 FILLER_0_48_370 ();
 FILLCELL_X1 FILLER_0_48_372 ();
 FILLCELL_X2 FILLER_0_48_383 ();
 FILLCELL_X2 FILLER_0_48_400 ();
 FILLCELL_X4 FILLER_0_48_436 ();
 FILLCELL_X4 FILLER_0_49_1 ();
 FILLCELL_X2 FILLER_0_49_15 ();
 FILLCELL_X1 FILLER_0_49_17 ();
 FILLCELL_X2 FILLER_0_49_61 ();
 FILLCELL_X1 FILLER_0_49_75 ();
 FILLCELL_X2 FILLER_0_49_94 ();
 FILLCELL_X4 FILLER_0_49_115 ();
 FILLCELL_X2 FILLER_0_49_119 ();
 FILLCELL_X2 FILLER_0_49_138 ();
 FILLCELL_X1 FILLER_0_49_144 ();
 FILLCELL_X2 FILLER_0_49_148 ();
 FILLCELL_X1 FILLER_0_49_150 ();
 FILLCELL_X1 FILLER_0_49_179 ();
 FILLCELL_X1 FILLER_0_49_183 ();
 FILLCELL_X2 FILLER_0_49_202 ();
 FILLCELL_X2 FILLER_0_49_208 ();
 FILLCELL_X1 FILLER_0_49_210 ();
 FILLCELL_X1 FILLER_0_49_218 ();
 FILLCELL_X1 FILLER_0_49_225 ();
 FILLCELL_X1 FILLER_0_49_229 ();
 FILLCELL_X2 FILLER_0_49_245 ();
 FILLCELL_X1 FILLER_0_49_247 ();
 FILLCELL_X1 FILLER_0_49_279 ();
 FILLCELL_X2 FILLER_0_49_286 ();
 FILLCELL_X1 FILLER_0_49_288 ();
 FILLCELL_X1 FILLER_0_49_294 ();
 FILLCELL_X1 FILLER_0_49_309 ();
 FILLCELL_X1 FILLER_0_49_313 ();
 FILLCELL_X1 FILLER_0_49_333 ();
 FILLCELL_X1 FILLER_0_49_344 ();
 FILLCELL_X8 FILLER_0_49_360 ();
 FILLCELL_X2 FILLER_0_49_368 ();
 FILLCELL_X1 FILLER_0_49_370 ();
 FILLCELL_X4 FILLER_0_49_379 ();
 FILLCELL_X1 FILLER_0_49_392 ();
 FILLCELL_X8 FILLER_0_49_400 ();
 FILLCELL_X4 FILLER_0_49_408 ();
 FILLCELL_X1 FILLER_0_49_412 ();
 FILLCELL_X2 FILLER_0_49_432 ();
 FILLCELL_X1 FILLER_0_50_1 ();
 FILLCELL_X1 FILLER_0_50_6 ();
 FILLCELL_X1 FILLER_0_50_17 ();
 FILLCELL_X2 FILLER_0_50_24 ();
 FILLCELL_X1 FILLER_0_50_26 ();
 FILLCELL_X2 FILLER_0_50_36 ();
 FILLCELL_X1 FILLER_0_50_54 ();
 FILLCELL_X4 FILLER_0_50_61 ();
 FILLCELL_X1 FILLER_0_50_71 ();
 FILLCELL_X2 FILLER_0_50_79 ();
 FILLCELL_X4 FILLER_0_50_85 ();
 FILLCELL_X8 FILLER_0_50_90 ();
 FILLCELL_X1 FILLER_0_50_98 ();
 FILLCELL_X4 FILLER_0_50_102 ();
 FILLCELL_X1 FILLER_0_50_106 ();
 FILLCELL_X16 FILLER_0_50_113 ();
 FILLCELL_X1 FILLER_0_50_146 ();
 FILLCELL_X2 FILLER_0_50_150 ();
 FILLCELL_X2 FILLER_0_50_201 ();
 FILLCELL_X1 FILLER_0_50_209 ();
 FILLCELL_X2 FILLER_0_50_227 ();
 FILLCELL_X1 FILLER_0_50_236 ();
 FILLCELL_X8 FILLER_0_50_247 ();
 FILLCELL_X4 FILLER_0_50_255 ();
 FILLCELL_X1 FILLER_0_50_259 ();
 FILLCELL_X4 FILLER_0_50_263 ();
 FILLCELL_X2 FILLER_0_50_284 ();
 FILLCELL_X2 FILLER_0_50_301 ();
 FILLCELL_X1 FILLER_0_50_310 ();
 FILLCELL_X4 FILLER_0_50_313 ();
 FILLCELL_X1 FILLER_0_50_317 ();
 FILLCELL_X2 FILLER_0_50_324 ();
 FILLCELL_X2 FILLER_0_50_329 ();
 FILLCELL_X1 FILLER_0_50_331 ();
 FILLCELL_X1 FILLER_0_50_341 ();
 FILLCELL_X1 FILLER_0_50_345 ();
 FILLCELL_X2 FILLER_0_50_369 ();
 FILLCELL_X1 FILLER_0_50_385 ();
 FILLCELL_X1 FILLER_0_50_389 ();
 FILLCELL_X4 FILLER_0_50_392 ();
 FILLCELL_X1 FILLER_0_50_396 ();
 FILLCELL_X8 FILLER_0_50_401 ();
 FILLCELL_X4 FILLER_0_50_409 ();
 FILLCELL_X2 FILLER_0_50_413 ();
 FILLCELL_X1 FILLER_0_50_415 ();
 FILLCELL_X1 FILLER_0_50_422 ();
 FILLCELL_X1 FILLER_0_51_1 ();
 FILLCELL_X1 FILLER_0_51_8 ();
 FILLCELL_X1 FILLER_0_51_18 ();
 FILLCELL_X2 FILLER_0_51_23 ();
 FILLCELL_X1 FILLER_0_51_25 ();
 FILLCELL_X2 FILLER_0_51_29 ();
 FILLCELL_X1 FILLER_0_51_31 ();
 FILLCELL_X2 FILLER_0_51_35 ();
 FILLCELL_X8 FILLER_0_51_47 ();
 FILLCELL_X1 FILLER_0_51_55 ();
 FILLCELL_X2 FILLER_0_51_86 ();
 FILLCELL_X2 FILLER_0_51_126 ();
 FILLCELL_X1 FILLER_0_51_130 ();
 FILLCELL_X1 FILLER_0_51_137 ();
 FILLCELL_X1 FILLER_0_51_141 ();
 FILLCELL_X8 FILLER_0_51_147 ();
 FILLCELL_X4 FILLER_0_51_155 ();
 FILLCELL_X2 FILLER_0_51_159 ();
 FILLCELL_X1 FILLER_0_51_166 ();
 FILLCELL_X1 FILLER_0_51_171 ();
 FILLCELL_X1 FILLER_0_51_179 ();
 FILLCELL_X1 FILLER_0_51_183 ();
 FILLCELL_X1 FILLER_0_51_190 ();
 FILLCELL_X1 FILLER_0_51_195 ();
 FILLCELL_X1 FILLER_0_51_201 ();
 FILLCELL_X1 FILLER_0_51_205 ();
 FILLCELL_X1 FILLER_0_51_209 ();
 FILLCELL_X2 FILLER_0_51_225 ();
 FILLCELL_X1 FILLER_0_51_236 ();
 FILLCELL_X1 FILLER_0_51_269 ();
 FILLCELL_X2 FILLER_0_51_283 ();
 FILLCELL_X1 FILLER_0_51_285 ();
 FILLCELL_X1 FILLER_0_51_292 ();
 FILLCELL_X1 FILLER_0_51_308 ();
 FILLCELL_X1 FILLER_0_51_345 ();
 FILLCELL_X4 FILLER_0_51_350 ();
 FILLCELL_X2 FILLER_0_51_354 ();
 FILLCELL_X1 FILLER_0_51_367 ();
 FILLCELL_X4 FILLER_0_51_385 ();
 FILLCELL_X1 FILLER_0_51_389 ();
 FILLCELL_X4 FILLER_0_51_410 ();
 FILLCELL_X2 FILLER_0_51_414 ();
 FILLCELL_X4 FILLER_0_52_1 ();
 FILLCELL_X2 FILLER_0_52_5 ();
 FILLCELL_X1 FILLER_0_52_7 ();
 FILLCELL_X1 FILLER_0_52_11 ();
 FILLCELL_X2 FILLER_0_52_16 ();
 FILLCELL_X2 FILLER_0_52_30 ();
 FILLCELL_X2 FILLER_0_52_50 ();
 FILLCELL_X1 FILLER_0_52_52 ();
 FILLCELL_X2 FILLER_0_52_87 ();
 FILLCELL_X1 FILLER_0_52_90 ();
 FILLCELL_X1 FILLER_0_52_97 ();
 FILLCELL_X1 FILLER_0_52_105 ();
 FILLCELL_X4 FILLER_0_52_112 ();
 FILLCELL_X1 FILLER_0_52_116 ();
 FILLCELL_X1 FILLER_0_52_144 ();
 FILLCELL_X8 FILLER_0_52_150 ();
 FILLCELL_X2 FILLER_0_52_158 ();
 FILLCELL_X2 FILLER_0_52_205 ();
 FILLCELL_X2 FILLER_0_52_211 ();
 FILLCELL_X1 FILLER_0_52_226 ();
 FILLCELL_X1 FILLER_0_52_231 ();
 FILLCELL_X1 FILLER_0_52_242 ();
 FILLCELL_X2 FILLER_0_52_250 ();
 FILLCELL_X1 FILLER_0_52_262 ();
 FILLCELL_X1 FILLER_0_52_266 ();
 FILLCELL_X2 FILLER_0_52_280 ();
 FILLCELL_X1 FILLER_0_52_285 ();
 FILLCELL_X4 FILLER_0_52_293 ();
 FILLCELL_X1 FILLER_0_52_297 ();
 FILLCELL_X1 FILLER_0_52_308 ();
 FILLCELL_X1 FILLER_0_52_313 ();
 FILLCELL_X2 FILLER_0_52_333 ();
 FILLCELL_X2 FILLER_0_52_344 ();
 FILLCELL_X1 FILLER_0_52_346 ();
 FILLCELL_X4 FILLER_0_52_351 ();
 FILLCELL_X2 FILLER_0_52_355 ();
 FILLCELL_X1 FILLER_0_52_357 ();
 FILLCELL_X2 FILLER_0_52_415 ();
 FILLCELL_X1 FILLER_0_52_417 ();
 FILLCELL_X1 FILLER_0_52_421 ();
 FILLCELL_X1 FILLER_0_52_439 ();
 FILLCELL_X2 FILLER_0_53_1 ();
 FILLCELL_X2 FILLER_0_53_30 ();
 FILLCELL_X1 FILLER_0_53_36 ();
 FILLCELL_X2 FILLER_0_53_43 ();
 FILLCELL_X2 FILLER_0_53_80 ();
 FILLCELL_X1 FILLER_0_53_82 ();
 FILLCELL_X8 FILLER_0_53_108 ();
 FILLCELL_X4 FILLER_0_53_147 ();
 FILLCELL_X2 FILLER_0_53_151 ();
 FILLCELL_X1 FILLER_0_53_153 ();
 FILLCELL_X4 FILLER_0_53_158 ();
 FILLCELL_X2 FILLER_0_53_232 ();
 FILLCELL_X1 FILLER_0_53_234 ();
 FILLCELL_X1 FILLER_0_53_258 ();
 FILLCELL_X2 FILLER_0_53_269 ();
 FILLCELL_X1 FILLER_0_53_290 ();
 FILLCELL_X2 FILLER_0_53_300 ();
 FILLCELL_X2 FILLER_0_53_308 ();
 FILLCELL_X4 FILLER_0_53_313 ();
 FILLCELL_X1 FILLER_0_53_317 ();
 FILLCELL_X2 FILLER_0_53_386 ();
 FILLCELL_X1 FILLER_0_53_388 ();
 FILLCELL_X1 FILLER_0_53_432 ();
 FILLCELL_X1 FILLER_0_53_436 ();
 FILLCELL_X4 FILLER_0_54_1 ();
 FILLCELL_X1 FILLER_0_54_5 ();
 FILLCELL_X1 FILLER_0_54_10 ();
 FILLCELL_X1 FILLER_0_54_15 ();
 FILLCELL_X1 FILLER_0_54_26 ();
 FILLCELL_X2 FILLER_0_54_58 ();
 FILLCELL_X1 FILLER_0_54_60 ();
 FILLCELL_X1 FILLER_0_54_83 ();
 FILLCELL_X8 FILLER_0_54_109 ();
 FILLCELL_X4 FILLER_0_54_117 ();
 FILLCELL_X4 FILLER_0_54_124 ();
 FILLCELL_X2 FILLER_0_54_128 ();
 FILLCELL_X4 FILLER_0_54_133 ();
 FILLCELL_X1 FILLER_0_54_143 ();
 FILLCELL_X2 FILLER_0_54_149 ();
 FILLCELL_X2 FILLER_0_54_154 ();
 FILLCELL_X2 FILLER_0_54_161 ();
 FILLCELL_X1 FILLER_0_54_163 ();
 FILLCELL_X1 FILLER_0_54_182 ();
 FILLCELL_X2 FILLER_0_54_192 ();
 FILLCELL_X2 FILLER_0_54_216 ();
 FILLCELL_X1 FILLER_0_54_225 ();
 FILLCELL_X4 FILLER_0_54_229 ();
 FILLCELL_X2 FILLER_0_54_261 ();
 FILLCELL_X1 FILLER_0_54_277 ();
 FILLCELL_X1 FILLER_0_54_284 ();
 FILLCELL_X1 FILLER_0_54_298 ();
 FILLCELL_X1 FILLER_0_54_310 ();
 FILLCELL_X1 FILLER_0_54_318 ();
 FILLCELL_X1 FILLER_0_54_322 ();
 FILLCELL_X1 FILLER_0_54_329 ();
 FILLCELL_X1 FILLER_0_54_350 ();
 FILLCELL_X1 FILLER_0_54_374 ();
 FILLCELL_X8 FILLER_0_54_382 ();
 FILLCELL_X2 FILLER_0_54_390 ();
 FILLCELL_X2 FILLER_0_54_434 ();
 FILLCELL_X16 FILLER_0_55_1 ();
 FILLCELL_X1 FILLER_0_55_17 ();
 FILLCELL_X8 FILLER_0_55_42 ();
 FILLCELL_X2 FILLER_0_55_93 ();
 FILLCELL_X2 FILLER_0_55_102 ();
 FILLCELL_X1 FILLER_0_55_104 ();
 FILLCELL_X1 FILLER_0_55_109 ();
 FILLCELL_X2 FILLER_0_55_119 ();
 FILLCELL_X1 FILLER_0_55_121 ();
 FILLCELL_X4 FILLER_0_55_149 ();
 FILLCELL_X8 FILLER_0_55_160 ();
 FILLCELL_X1 FILLER_0_55_168 ();
 FILLCELL_X2 FILLER_0_55_175 ();
 FILLCELL_X1 FILLER_0_55_177 ();
 FILLCELL_X4 FILLER_0_55_179 ();
 FILLCELL_X2 FILLER_0_55_189 ();
 FILLCELL_X1 FILLER_0_55_191 ();
 FILLCELL_X1 FILLER_0_55_195 ();
 FILLCELL_X1 FILLER_0_55_200 ();
 FILLCELL_X1 FILLER_0_55_207 ();
 FILLCELL_X1 FILLER_0_55_211 ();
 FILLCELL_X2 FILLER_0_55_225 ();
 FILLCELL_X1 FILLER_0_55_227 ();
 FILLCELL_X1 FILLER_0_55_237 ();
 FILLCELL_X1 FILLER_0_55_244 ();
 FILLCELL_X1 FILLER_0_55_248 ();
 FILLCELL_X1 FILLER_0_55_255 ();
 FILLCELL_X1 FILLER_0_55_259 ();
 FILLCELL_X4 FILLER_0_55_266 ();
 FILLCELL_X1 FILLER_0_55_270 ();
 FILLCELL_X1 FILLER_0_55_280 ();
 FILLCELL_X1 FILLER_0_55_285 ();
 FILLCELL_X1 FILLER_0_55_295 ();
 FILLCELL_X1 FILLER_0_55_299 ();
 FILLCELL_X1 FILLER_0_55_306 ();
 FILLCELL_X1 FILLER_0_55_310 ();
 FILLCELL_X1 FILLER_0_55_320 ();
 FILLCELL_X1 FILLER_0_55_330 ();
 FILLCELL_X2 FILLER_0_55_337 ();
 FILLCELL_X1 FILLER_0_55_345 ();
 FILLCELL_X1 FILLER_0_55_364 ();
 FILLCELL_X1 FILLER_0_55_369 ();
 FILLCELL_X1 FILLER_0_55_390 ();
 FILLCELL_X1 FILLER_0_55_394 ();
 FILLCELL_X1 FILLER_0_55_399 ();
 FILLCELL_X1 FILLER_0_55_403 ();
 FILLCELL_X1 FILLER_0_55_408 ();
 FILLCELL_X2 FILLER_0_55_412 ();
 FILLCELL_X1 FILLER_0_55_417 ();
 FILLCELL_X2 FILLER_0_55_421 ();
 FILLCELL_X1 FILLER_0_56_1 ();
 FILLCELL_X4 FILLER_0_56_19 ();
 FILLCELL_X2 FILLER_0_56_36 ();
 FILLCELL_X1 FILLER_0_56_38 ();
 FILLCELL_X8 FILLER_0_56_43 ();
 FILLCELL_X4 FILLER_0_56_51 ();
 FILLCELL_X2 FILLER_0_56_55 ();
 FILLCELL_X2 FILLER_0_56_60 ();
 FILLCELL_X1 FILLER_0_56_62 ();
 FILLCELL_X1 FILLER_0_56_88 ();
 FILLCELL_X2 FILLER_0_56_93 ();
 FILLCELL_X2 FILLER_0_56_107 ();
 FILLCELL_X1 FILLER_0_56_109 ();
 FILLCELL_X2 FILLER_0_56_137 ();
 FILLCELL_X16 FILLER_0_56_153 ();
 FILLCELL_X4 FILLER_0_56_169 ();
 FILLCELL_X1 FILLER_0_56_173 ();
 FILLCELL_X4 FILLER_0_56_214 ();
 FILLCELL_X2 FILLER_0_56_218 ();
 FILLCELL_X1 FILLER_0_56_223 ();
 FILLCELL_X2 FILLER_0_56_241 ();
 FILLCELL_X2 FILLER_0_56_273 ();
 FILLCELL_X2 FILLER_0_56_278 ();
 FILLCELL_X1 FILLER_0_56_286 ();
 FILLCELL_X4 FILLER_0_56_293 ();
 FILLCELL_X1 FILLER_0_56_297 ();
 FILLCELL_X1 FILLER_0_56_312 ();
 FILLCELL_X1 FILLER_0_56_327 ();
 FILLCELL_X2 FILLER_0_56_361 ();
 FILLCELL_X1 FILLER_0_56_363 ();
 FILLCELL_X1 FILLER_0_56_377 ();
 FILLCELL_X2 FILLER_0_56_381 ();
 FILLCELL_X1 FILLER_0_56_386 ();
 FILLCELL_X2 FILLER_0_56_404 ();
 FILLCELL_X2 FILLER_0_56_409 ();
 FILLCELL_X2 FILLER_0_56_415 ();
 FILLCELL_X2 FILLER_0_56_420 ();
 FILLCELL_X1 FILLER_0_56_422 ();
 FILLCELL_X4 FILLER_0_56_429 ();
 FILLCELL_X1 FILLER_0_56_433 ();
 FILLCELL_X16 FILLER_0_57_1 ();
 FILLCELL_X4 FILLER_0_57_17 ();
 FILLCELL_X2 FILLER_0_57_21 ();
 FILLCELL_X1 FILLER_0_57_23 ();
 FILLCELL_X16 FILLER_0_57_44 ();
 FILLCELL_X8 FILLER_0_57_60 ();
 FILLCELL_X4 FILLER_0_57_68 ();
 FILLCELL_X1 FILLER_0_57_72 ();
 FILLCELL_X2 FILLER_0_57_76 ();
 FILLCELL_X1 FILLER_0_57_95 ();
 FILLCELL_X1 FILLER_0_57_99 ();
 FILLCELL_X8 FILLER_0_57_106 ();
 FILLCELL_X1 FILLER_0_57_114 ();
 FILLCELL_X1 FILLER_0_57_121 ();
 FILLCELL_X16 FILLER_0_57_125 ();
 FILLCELL_X2 FILLER_0_57_141 ();
 FILLCELL_X1 FILLER_0_57_143 ();
 FILLCELL_X16 FILLER_0_57_161 ();
 FILLCELL_X1 FILLER_0_57_177 ();
 FILLCELL_X1 FILLER_0_57_179 ();
 FILLCELL_X8 FILLER_0_57_197 ();
 FILLCELL_X2 FILLER_0_57_205 ();
 FILLCELL_X1 FILLER_0_57_224 ();
 FILLCELL_X2 FILLER_0_57_230 ();
 FILLCELL_X1 FILLER_0_57_238 ();
 FILLCELL_X1 FILLER_0_57_242 ();
 FILLCELL_X2 FILLER_0_57_272 ();
 FILLCELL_X1 FILLER_0_57_302 ();
 FILLCELL_X4 FILLER_0_57_345 ();
 FILLCELL_X1 FILLER_0_57_349 ();
 FILLCELL_X1 FILLER_0_57_359 ();
 FILLCELL_X1 FILLER_0_57_377 ();
 FILLCELL_X2 FILLER_0_57_402 ();
 FILLCELL_X1 FILLER_0_57_404 ();
 FILLCELL_X2 FILLER_0_57_422 ();
 FILLCELL_X8 FILLER_0_57_431 ();
 FILLCELL_X1 FILLER_0_57_439 ();
 FILLCELL_X32 FILLER_0_58_1 ();
 FILLCELL_X4 FILLER_0_58_33 ();
 FILLCELL_X2 FILLER_0_58_37 ();
 FILLCELL_X16 FILLER_0_58_56 ();
 FILLCELL_X4 FILLER_0_58_72 ();
 FILLCELL_X1 FILLER_0_58_76 ();
 FILLCELL_X2 FILLER_0_58_86 ();
 FILLCELL_X1 FILLER_0_58_88 ();
 FILLCELL_X4 FILLER_0_58_90 ();
 FILLCELL_X2 FILLER_0_58_94 ();
 FILLCELL_X32 FILLER_0_58_108 ();
 FILLCELL_X16 FILLER_0_58_140 ();
 FILLCELL_X4 FILLER_0_58_156 ();
 FILLCELL_X2 FILLER_0_58_166 ();
 FILLCELL_X4 FILLER_0_58_171 ();
 FILLCELL_X2 FILLER_0_58_175 ();
 FILLCELL_X1 FILLER_0_58_177 ();
 FILLCELL_X8 FILLER_0_58_179 ();
 FILLCELL_X2 FILLER_0_58_187 ();
 FILLCELL_X1 FILLER_0_58_189 ();
 FILLCELL_X4 FILLER_0_58_193 ();
 FILLCELL_X1 FILLER_0_58_197 ();
 FILLCELL_X1 FILLER_0_58_213 ();
 FILLCELL_X4 FILLER_0_58_233 ();
 FILLCELL_X1 FILLER_0_58_237 ();
 FILLCELL_X2 FILLER_0_58_241 ();
 FILLCELL_X1 FILLER_0_58_243 ();
 FILLCELL_X4 FILLER_0_58_271 ();
 FILLCELL_X2 FILLER_0_58_321 ();
 FILLCELL_X1 FILLER_0_58_323 ();
 FILLCELL_X2 FILLER_0_58_330 ();
 FILLCELL_X1 FILLER_0_58_340 ();
 FILLCELL_X1 FILLER_0_58_345 ();
 FILLCELL_X1 FILLER_0_58_355 ();
 FILLCELL_X8 FILLER_0_58_357 ();
 FILLCELL_X8 FILLER_0_58_405 ();
 FILLCELL_X2 FILLER_0_58_413 ();
 FILLCELL_X1 FILLER_0_58_415 ();
 FILLCELL_X4 FILLER_0_58_433 ();
 FILLCELL_X2 FILLER_0_58_437 ();
 FILLCELL_X1 FILLER_0_58_439 ();
endmodule
